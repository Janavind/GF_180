magic
tech gf180mcuC
magscale 1 5
timestamp 1670269577
<< obsm1 >>
rect 672 855 59304 58617
<< metal2 >>
rect 1232 59600 1288 60000
rect 1736 59600 1792 60000
rect 2240 59600 2296 60000
rect 2744 59600 2800 60000
rect 3248 59600 3304 60000
rect 3752 59600 3808 60000
rect 4256 59600 4312 60000
rect 4760 59600 4816 60000
rect 5264 59600 5320 60000
rect 5768 59600 5824 60000
rect 6272 59600 6328 60000
rect 6776 59600 6832 60000
rect 7280 59600 7336 60000
rect 7784 59600 7840 60000
rect 8288 59600 8344 60000
rect 8792 59600 8848 60000
rect 9296 59600 9352 60000
rect 9800 59600 9856 60000
rect 10304 59600 10360 60000
rect 10808 59600 10864 60000
rect 11312 59600 11368 60000
rect 11816 59600 11872 60000
rect 12320 59600 12376 60000
rect 12824 59600 12880 60000
rect 13328 59600 13384 60000
rect 13832 59600 13888 60000
rect 14336 59600 14392 60000
rect 14840 59600 14896 60000
rect 15344 59600 15400 60000
rect 15848 59600 15904 60000
rect 16352 59600 16408 60000
rect 16856 59600 16912 60000
rect 17360 59600 17416 60000
rect 17864 59600 17920 60000
rect 18368 59600 18424 60000
rect 18872 59600 18928 60000
rect 19376 59600 19432 60000
rect 19880 59600 19936 60000
rect 20384 59600 20440 60000
rect 20888 59600 20944 60000
rect 21392 59600 21448 60000
rect 21896 59600 21952 60000
rect 22400 59600 22456 60000
rect 22904 59600 22960 60000
rect 23408 59600 23464 60000
rect 23912 59600 23968 60000
rect 24416 59600 24472 60000
rect 24920 59600 24976 60000
rect 25424 59600 25480 60000
rect 25928 59600 25984 60000
rect 26432 59600 26488 60000
rect 26936 59600 26992 60000
rect 27440 59600 27496 60000
rect 27944 59600 28000 60000
rect 28448 59600 28504 60000
rect 28952 59600 29008 60000
rect 29456 59600 29512 60000
rect 29960 59600 30016 60000
rect 30464 59600 30520 60000
rect 30968 59600 31024 60000
rect 31472 59600 31528 60000
rect 31976 59600 32032 60000
rect 32480 59600 32536 60000
rect 32984 59600 33040 60000
rect 33488 59600 33544 60000
rect 33992 59600 34048 60000
rect 34496 59600 34552 60000
rect 35000 59600 35056 60000
rect 35504 59600 35560 60000
rect 36008 59600 36064 60000
rect 36512 59600 36568 60000
rect 37016 59600 37072 60000
rect 37520 59600 37576 60000
rect 38024 59600 38080 60000
rect 38528 59600 38584 60000
rect 39032 59600 39088 60000
rect 39536 59600 39592 60000
rect 40040 59600 40096 60000
rect 40544 59600 40600 60000
rect 41048 59600 41104 60000
rect 41552 59600 41608 60000
rect 42056 59600 42112 60000
rect 42560 59600 42616 60000
rect 43064 59600 43120 60000
rect 43568 59600 43624 60000
rect 44072 59600 44128 60000
rect 44576 59600 44632 60000
rect 45080 59600 45136 60000
rect 45584 59600 45640 60000
rect 46088 59600 46144 60000
rect 46592 59600 46648 60000
rect 47096 59600 47152 60000
rect 47600 59600 47656 60000
rect 48104 59600 48160 60000
rect 48608 59600 48664 60000
rect 49112 59600 49168 60000
rect 49616 59600 49672 60000
rect 50120 59600 50176 60000
rect 50624 59600 50680 60000
rect 51128 59600 51184 60000
rect 51632 59600 51688 60000
rect 52136 59600 52192 60000
rect 52640 59600 52696 60000
rect 53144 59600 53200 60000
rect 53648 59600 53704 60000
rect 54152 59600 54208 60000
rect 54656 59600 54712 60000
rect 55160 59600 55216 60000
rect 55664 59600 55720 60000
rect 56168 59600 56224 60000
rect 56672 59600 56728 60000
rect 57176 59600 57232 60000
rect 57680 59600 57736 60000
rect 58184 59600 58240 60000
rect 58688 59600 58744 60000
rect 4760 0 4816 400
rect 4928 0 4984 400
rect 5096 0 5152 400
rect 5264 0 5320 400
rect 5432 0 5488 400
rect 5600 0 5656 400
rect 5768 0 5824 400
rect 5936 0 5992 400
rect 6104 0 6160 400
rect 6272 0 6328 400
rect 6440 0 6496 400
rect 6608 0 6664 400
rect 6776 0 6832 400
rect 6944 0 7000 400
rect 7112 0 7168 400
rect 7280 0 7336 400
rect 7448 0 7504 400
rect 7616 0 7672 400
rect 7784 0 7840 400
rect 7952 0 8008 400
rect 8120 0 8176 400
rect 8288 0 8344 400
rect 8456 0 8512 400
rect 8624 0 8680 400
rect 8792 0 8848 400
rect 8960 0 9016 400
rect 9128 0 9184 400
rect 9296 0 9352 400
rect 9464 0 9520 400
rect 9632 0 9688 400
rect 9800 0 9856 400
rect 9968 0 10024 400
rect 10136 0 10192 400
rect 10304 0 10360 400
rect 10472 0 10528 400
rect 10640 0 10696 400
rect 10808 0 10864 400
rect 10976 0 11032 400
rect 11144 0 11200 400
rect 11312 0 11368 400
rect 11480 0 11536 400
rect 11648 0 11704 400
rect 11816 0 11872 400
rect 11984 0 12040 400
rect 12152 0 12208 400
rect 12320 0 12376 400
rect 12488 0 12544 400
rect 12656 0 12712 400
rect 12824 0 12880 400
rect 12992 0 13048 400
rect 13160 0 13216 400
rect 13328 0 13384 400
rect 13496 0 13552 400
rect 13664 0 13720 400
rect 13832 0 13888 400
rect 14000 0 14056 400
rect 14168 0 14224 400
rect 14336 0 14392 400
rect 14504 0 14560 400
rect 14672 0 14728 400
rect 14840 0 14896 400
rect 15008 0 15064 400
rect 15176 0 15232 400
rect 15344 0 15400 400
rect 15512 0 15568 400
rect 15680 0 15736 400
rect 15848 0 15904 400
rect 16016 0 16072 400
rect 16184 0 16240 400
rect 16352 0 16408 400
rect 16520 0 16576 400
rect 16688 0 16744 400
rect 16856 0 16912 400
rect 17024 0 17080 400
rect 17192 0 17248 400
rect 17360 0 17416 400
rect 17528 0 17584 400
rect 17696 0 17752 400
rect 17864 0 17920 400
rect 18032 0 18088 400
rect 18200 0 18256 400
rect 18368 0 18424 400
rect 18536 0 18592 400
rect 18704 0 18760 400
rect 18872 0 18928 400
rect 19040 0 19096 400
rect 19208 0 19264 400
rect 19376 0 19432 400
rect 19544 0 19600 400
rect 19712 0 19768 400
rect 19880 0 19936 400
rect 20048 0 20104 400
rect 20216 0 20272 400
rect 20384 0 20440 400
rect 20552 0 20608 400
rect 20720 0 20776 400
rect 20888 0 20944 400
rect 21056 0 21112 400
rect 21224 0 21280 400
rect 21392 0 21448 400
rect 21560 0 21616 400
rect 21728 0 21784 400
rect 21896 0 21952 400
rect 22064 0 22120 400
rect 22232 0 22288 400
rect 22400 0 22456 400
rect 22568 0 22624 400
rect 22736 0 22792 400
rect 22904 0 22960 400
rect 23072 0 23128 400
rect 23240 0 23296 400
rect 23408 0 23464 400
rect 23576 0 23632 400
rect 23744 0 23800 400
rect 23912 0 23968 400
rect 24080 0 24136 400
rect 24248 0 24304 400
rect 24416 0 24472 400
rect 24584 0 24640 400
rect 24752 0 24808 400
rect 24920 0 24976 400
rect 25088 0 25144 400
rect 25256 0 25312 400
rect 25424 0 25480 400
rect 25592 0 25648 400
rect 25760 0 25816 400
rect 25928 0 25984 400
rect 26096 0 26152 400
rect 26264 0 26320 400
rect 26432 0 26488 400
rect 26600 0 26656 400
rect 26768 0 26824 400
rect 26936 0 26992 400
rect 27104 0 27160 400
rect 27272 0 27328 400
rect 27440 0 27496 400
rect 27608 0 27664 400
rect 27776 0 27832 400
rect 27944 0 28000 400
rect 28112 0 28168 400
rect 28280 0 28336 400
rect 28448 0 28504 400
rect 28616 0 28672 400
rect 28784 0 28840 400
rect 28952 0 29008 400
rect 29120 0 29176 400
rect 29288 0 29344 400
rect 29456 0 29512 400
rect 29624 0 29680 400
rect 29792 0 29848 400
rect 29960 0 30016 400
rect 30128 0 30184 400
rect 30296 0 30352 400
rect 30464 0 30520 400
rect 30632 0 30688 400
rect 30800 0 30856 400
rect 30968 0 31024 400
rect 31136 0 31192 400
rect 31304 0 31360 400
rect 31472 0 31528 400
rect 31640 0 31696 400
rect 31808 0 31864 400
rect 31976 0 32032 400
rect 32144 0 32200 400
rect 32312 0 32368 400
rect 32480 0 32536 400
rect 32648 0 32704 400
rect 32816 0 32872 400
rect 32984 0 33040 400
rect 33152 0 33208 400
rect 33320 0 33376 400
rect 33488 0 33544 400
rect 33656 0 33712 400
rect 33824 0 33880 400
rect 33992 0 34048 400
rect 34160 0 34216 400
rect 34328 0 34384 400
rect 34496 0 34552 400
rect 34664 0 34720 400
rect 34832 0 34888 400
rect 35000 0 35056 400
rect 35168 0 35224 400
rect 35336 0 35392 400
rect 35504 0 35560 400
rect 35672 0 35728 400
rect 35840 0 35896 400
rect 36008 0 36064 400
rect 36176 0 36232 400
rect 36344 0 36400 400
rect 36512 0 36568 400
rect 36680 0 36736 400
rect 36848 0 36904 400
rect 37016 0 37072 400
rect 37184 0 37240 400
rect 37352 0 37408 400
rect 37520 0 37576 400
rect 37688 0 37744 400
rect 37856 0 37912 400
rect 38024 0 38080 400
rect 38192 0 38248 400
rect 38360 0 38416 400
rect 38528 0 38584 400
rect 38696 0 38752 400
rect 38864 0 38920 400
rect 39032 0 39088 400
rect 39200 0 39256 400
rect 39368 0 39424 400
rect 39536 0 39592 400
rect 39704 0 39760 400
rect 39872 0 39928 400
rect 40040 0 40096 400
rect 40208 0 40264 400
rect 40376 0 40432 400
rect 40544 0 40600 400
rect 40712 0 40768 400
rect 40880 0 40936 400
rect 41048 0 41104 400
rect 41216 0 41272 400
rect 41384 0 41440 400
rect 41552 0 41608 400
rect 41720 0 41776 400
rect 41888 0 41944 400
rect 42056 0 42112 400
rect 42224 0 42280 400
rect 42392 0 42448 400
rect 42560 0 42616 400
rect 42728 0 42784 400
rect 42896 0 42952 400
rect 43064 0 43120 400
rect 43232 0 43288 400
rect 43400 0 43456 400
rect 43568 0 43624 400
rect 43736 0 43792 400
rect 43904 0 43960 400
rect 44072 0 44128 400
rect 44240 0 44296 400
rect 44408 0 44464 400
rect 44576 0 44632 400
rect 44744 0 44800 400
rect 44912 0 44968 400
rect 45080 0 45136 400
rect 45248 0 45304 400
rect 45416 0 45472 400
rect 45584 0 45640 400
rect 45752 0 45808 400
rect 45920 0 45976 400
rect 46088 0 46144 400
rect 46256 0 46312 400
rect 46424 0 46480 400
rect 46592 0 46648 400
rect 46760 0 46816 400
rect 46928 0 46984 400
rect 47096 0 47152 400
rect 47264 0 47320 400
rect 47432 0 47488 400
rect 47600 0 47656 400
rect 47768 0 47824 400
rect 47936 0 47992 400
rect 48104 0 48160 400
rect 48272 0 48328 400
rect 48440 0 48496 400
rect 48608 0 48664 400
rect 48776 0 48832 400
rect 48944 0 49000 400
rect 49112 0 49168 400
rect 49280 0 49336 400
rect 49448 0 49504 400
rect 49616 0 49672 400
rect 49784 0 49840 400
rect 49952 0 50008 400
rect 50120 0 50176 400
rect 50288 0 50344 400
rect 50456 0 50512 400
rect 50624 0 50680 400
rect 50792 0 50848 400
rect 50960 0 51016 400
rect 51128 0 51184 400
rect 51296 0 51352 400
rect 51464 0 51520 400
rect 51632 0 51688 400
rect 51800 0 51856 400
rect 51968 0 52024 400
rect 52136 0 52192 400
rect 52304 0 52360 400
rect 52472 0 52528 400
rect 52640 0 52696 400
rect 52808 0 52864 400
rect 52976 0 53032 400
rect 53144 0 53200 400
rect 53312 0 53368 400
rect 53480 0 53536 400
rect 53648 0 53704 400
rect 53816 0 53872 400
rect 53984 0 54040 400
rect 54152 0 54208 400
rect 54320 0 54376 400
rect 54488 0 54544 400
rect 54656 0 54712 400
rect 54824 0 54880 400
rect 54992 0 55048 400
rect 55160 0 55216 400
<< obsm2 >>
rect 2326 59570 2714 59600
rect 2830 59570 3218 59600
rect 3334 59570 3722 59600
rect 3838 59570 4226 59600
rect 4342 59570 4730 59600
rect 4846 59570 5234 59600
rect 5350 59570 5738 59600
rect 5854 59570 6242 59600
rect 6358 59570 6746 59600
rect 6862 59570 7250 59600
rect 7366 59570 7754 59600
rect 7870 59570 8258 59600
rect 8374 59570 8762 59600
rect 8878 59570 9266 59600
rect 9382 59570 9770 59600
rect 9886 59570 10274 59600
rect 10390 59570 10778 59600
rect 10894 59570 11282 59600
rect 11398 59570 11786 59600
rect 11902 59570 12290 59600
rect 12406 59570 12794 59600
rect 12910 59570 13298 59600
rect 13414 59570 13802 59600
rect 13918 59570 14306 59600
rect 14422 59570 14810 59600
rect 14926 59570 15314 59600
rect 15430 59570 15818 59600
rect 15934 59570 16322 59600
rect 16438 59570 16826 59600
rect 16942 59570 17330 59600
rect 17446 59570 17834 59600
rect 17950 59570 18338 59600
rect 18454 59570 18842 59600
rect 18958 59570 19346 59600
rect 19462 59570 19850 59600
rect 19966 59570 20354 59600
rect 20470 59570 20858 59600
rect 20974 59570 21362 59600
rect 21478 59570 21866 59600
rect 21982 59570 22370 59600
rect 22486 59570 22874 59600
rect 22990 59570 23378 59600
rect 23494 59570 23882 59600
rect 23998 59570 24386 59600
rect 24502 59570 24890 59600
rect 25006 59570 25394 59600
rect 25510 59570 25898 59600
rect 26014 59570 26402 59600
rect 26518 59570 26906 59600
rect 27022 59570 27410 59600
rect 27526 59570 27914 59600
rect 28030 59570 28418 59600
rect 28534 59570 28922 59600
rect 29038 59570 29426 59600
rect 29542 59570 29930 59600
rect 30046 59570 30434 59600
rect 30550 59570 30938 59600
rect 31054 59570 31442 59600
rect 31558 59570 31946 59600
rect 32062 59570 32450 59600
rect 32566 59570 32954 59600
rect 33070 59570 33458 59600
rect 33574 59570 33962 59600
rect 34078 59570 34466 59600
rect 34582 59570 34970 59600
rect 35086 59570 35474 59600
rect 35590 59570 35978 59600
rect 36094 59570 36482 59600
rect 36598 59570 36986 59600
rect 37102 59570 37490 59600
rect 37606 59570 37994 59600
rect 38110 59570 38498 59600
rect 38614 59570 39002 59600
rect 39118 59570 39506 59600
rect 39622 59570 40010 59600
rect 40126 59570 40514 59600
rect 40630 59570 41018 59600
rect 41134 59570 41522 59600
rect 41638 59570 42026 59600
rect 42142 59570 42530 59600
rect 42646 59570 43034 59600
rect 43150 59570 43538 59600
rect 43654 59570 44042 59600
rect 44158 59570 44546 59600
rect 44662 59570 45050 59600
rect 45166 59570 45554 59600
rect 45670 59570 46058 59600
rect 46174 59570 46562 59600
rect 46678 59570 47066 59600
rect 47182 59570 47570 59600
rect 47686 59570 48074 59600
rect 48190 59570 48578 59600
rect 48694 59570 49082 59600
rect 49198 59570 49586 59600
rect 49702 59570 50090 59600
rect 50206 59570 50594 59600
rect 50710 59570 51098 59600
rect 51214 59570 51602 59600
rect 51718 59570 52106 59600
rect 52222 59570 52610 59600
rect 52726 59570 53114 59600
rect 53230 59570 53618 59600
rect 53734 59570 54122 59600
rect 54238 59570 54626 59600
rect 54742 59570 55130 59600
rect 55246 59570 55634 59600
rect 55750 59570 56138 59600
rect 56254 59570 56642 59600
rect 56758 59570 57146 59600
rect 57262 59570 57650 59600
rect 57766 59570 58154 59600
rect 58270 59570 58658 59600
rect 58774 59570 58842 59600
rect 2238 430 58842 59570
rect 2238 400 4730 430
rect 4846 400 4898 430
rect 5014 400 5066 430
rect 5182 400 5234 430
rect 5350 400 5402 430
rect 5518 400 5570 430
rect 5686 400 5738 430
rect 5854 400 5906 430
rect 6022 400 6074 430
rect 6190 400 6242 430
rect 6358 400 6410 430
rect 6526 400 6578 430
rect 6694 400 6746 430
rect 6862 400 6914 430
rect 7030 400 7082 430
rect 7198 400 7250 430
rect 7366 400 7418 430
rect 7534 400 7586 430
rect 7702 400 7754 430
rect 7870 400 7922 430
rect 8038 400 8090 430
rect 8206 400 8258 430
rect 8374 400 8426 430
rect 8542 400 8594 430
rect 8710 400 8762 430
rect 8878 400 8930 430
rect 9046 400 9098 430
rect 9214 400 9266 430
rect 9382 400 9434 430
rect 9550 400 9602 430
rect 9718 400 9770 430
rect 9886 400 9938 430
rect 10054 400 10106 430
rect 10222 400 10274 430
rect 10390 400 10442 430
rect 10558 400 10610 430
rect 10726 400 10778 430
rect 10894 400 10946 430
rect 11062 400 11114 430
rect 11230 400 11282 430
rect 11398 400 11450 430
rect 11566 400 11618 430
rect 11734 400 11786 430
rect 11902 400 11954 430
rect 12070 400 12122 430
rect 12238 400 12290 430
rect 12406 400 12458 430
rect 12574 400 12626 430
rect 12742 400 12794 430
rect 12910 400 12962 430
rect 13078 400 13130 430
rect 13246 400 13298 430
rect 13414 400 13466 430
rect 13582 400 13634 430
rect 13750 400 13802 430
rect 13918 400 13970 430
rect 14086 400 14138 430
rect 14254 400 14306 430
rect 14422 400 14474 430
rect 14590 400 14642 430
rect 14758 400 14810 430
rect 14926 400 14978 430
rect 15094 400 15146 430
rect 15262 400 15314 430
rect 15430 400 15482 430
rect 15598 400 15650 430
rect 15766 400 15818 430
rect 15934 400 15986 430
rect 16102 400 16154 430
rect 16270 400 16322 430
rect 16438 400 16490 430
rect 16606 400 16658 430
rect 16774 400 16826 430
rect 16942 400 16994 430
rect 17110 400 17162 430
rect 17278 400 17330 430
rect 17446 400 17498 430
rect 17614 400 17666 430
rect 17782 400 17834 430
rect 17950 400 18002 430
rect 18118 400 18170 430
rect 18286 400 18338 430
rect 18454 400 18506 430
rect 18622 400 18674 430
rect 18790 400 18842 430
rect 18958 400 19010 430
rect 19126 400 19178 430
rect 19294 400 19346 430
rect 19462 400 19514 430
rect 19630 400 19682 430
rect 19798 400 19850 430
rect 19966 400 20018 430
rect 20134 400 20186 430
rect 20302 400 20354 430
rect 20470 400 20522 430
rect 20638 400 20690 430
rect 20806 400 20858 430
rect 20974 400 21026 430
rect 21142 400 21194 430
rect 21310 400 21362 430
rect 21478 400 21530 430
rect 21646 400 21698 430
rect 21814 400 21866 430
rect 21982 400 22034 430
rect 22150 400 22202 430
rect 22318 400 22370 430
rect 22486 400 22538 430
rect 22654 400 22706 430
rect 22822 400 22874 430
rect 22990 400 23042 430
rect 23158 400 23210 430
rect 23326 400 23378 430
rect 23494 400 23546 430
rect 23662 400 23714 430
rect 23830 400 23882 430
rect 23998 400 24050 430
rect 24166 400 24218 430
rect 24334 400 24386 430
rect 24502 400 24554 430
rect 24670 400 24722 430
rect 24838 400 24890 430
rect 25006 400 25058 430
rect 25174 400 25226 430
rect 25342 400 25394 430
rect 25510 400 25562 430
rect 25678 400 25730 430
rect 25846 400 25898 430
rect 26014 400 26066 430
rect 26182 400 26234 430
rect 26350 400 26402 430
rect 26518 400 26570 430
rect 26686 400 26738 430
rect 26854 400 26906 430
rect 27022 400 27074 430
rect 27190 400 27242 430
rect 27358 400 27410 430
rect 27526 400 27578 430
rect 27694 400 27746 430
rect 27862 400 27914 430
rect 28030 400 28082 430
rect 28198 400 28250 430
rect 28366 400 28418 430
rect 28534 400 28586 430
rect 28702 400 28754 430
rect 28870 400 28922 430
rect 29038 400 29090 430
rect 29206 400 29258 430
rect 29374 400 29426 430
rect 29542 400 29594 430
rect 29710 400 29762 430
rect 29878 400 29930 430
rect 30046 400 30098 430
rect 30214 400 30266 430
rect 30382 400 30434 430
rect 30550 400 30602 430
rect 30718 400 30770 430
rect 30886 400 30938 430
rect 31054 400 31106 430
rect 31222 400 31274 430
rect 31390 400 31442 430
rect 31558 400 31610 430
rect 31726 400 31778 430
rect 31894 400 31946 430
rect 32062 400 32114 430
rect 32230 400 32282 430
rect 32398 400 32450 430
rect 32566 400 32618 430
rect 32734 400 32786 430
rect 32902 400 32954 430
rect 33070 400 33122 430
rect 33238 400 33290 430
rect 33406 400 33458 430
rect 33574 400 33626 430
rect 33742 400 33794 430
rect 33910 400 33962 430
rect 34078 400 34130 430
rect 34246 400 34298 430
rect 34414 400 34466 430
rect 34582 400 34634 430
rect 34750 400 34802 430
rect 34918 400 34970 430
rect 35086 400 35138 430
rect 35254 400 35306 430
rect 35422 400 35474 430
rect 35590 400 35642 430
rect 35758 400 35810 430
rect 35926 400 35978 430
rect 36094 400 36146 430
rect 36262 400 36314 430
rect 36430 400 36482 430
rect 36598 400 36650 430
rect 36766 400 36818 430
rect 36934 400 36986 430
rect 37102 400 37154 430
rect 37270 400 37322 430
rect 37438 400 37490 430
rect 37606 400 37658 430
rect 37774 400 37826 430
rect 37942 400 37994 430
rect 38110 400 38162 430
rect 38278 400 38330 430
rect 38446 400 38498 430
rect 38614 400 38666 430
rect 38782 400 38834 430
rect 38950 400 39002 430
rect 39118 400 39170 430
rect 39286 400 39338 430
rect 39454 400 39506 430
rect 39622 400 39674 430
rect 39790 400 39842 430
rect 39958 400 40010 430
rect 40126 400 40178 430
rect 40294 400 40346 430
rect 40462 400 40514 430
rect 40630 400 40682 430
rect 40798 400 40850 430
rect 40966 400 41018 430
rect 41134 400 41186 430
rect 41302 400 41354 430
rect 41470 400 41522 430
rect 41638 400 41690 430
rect 41806 400 41858 430
rect 41974 400 42026 430
rect 42142 400 42194 430
rect 42310 400 42362 430
rect 42478 400 42530 430
rect 42646 400 42698 430
rect 42814 400 42866 430
rect 42982 400 43034 430
rect 43150 400 43202 430
rect 43318 400 43370 430
rect 43486 400 43538 430
rect 43654 400 43706 430
rect 43822 400 43874 430
rect 43990 400 44042 430
rect 44158 400 44210 430
rect 44326 400 44378 430
rect 44494 400 44546 430
rect 44662 400 44714 430
rect 44830 400 44882 430
rect 44998 400 45050 430
rect 45166 400 45218 430
rect 45334 400 45386 430
rect 45502 400 45554 430
rect 45670 400 45722 430
rect 45838 400 45890 430
rect 46006 400 46058 430
rect 46174 400 46226 430
rect 46342 400 46394 430
rect 46510 400 46562 430
rect 46678 400 46730 430
rect 46846 400 46898 430
rect 47014 400 47066 430
rect 47182 400 47234 430
rect 47350 400 47402 430
rect 47518 400 47570 430
rect 47686 400 47738 430
rect 47854 400 47906 430
rect 48022 400 48074 430
rect 48190 400 48242 430
rect 48358 400 48410 430
rect 48526 400 48578 430
rect 48694 400 48746 430
rect 48862 400 48914 430
rect 49030 400 49082 430
rect 49198 400 49250 430
rect 49366 400 49418 430
rect 49534 400 49586 430
rect 49702 400 49754 430
rect 49870 400 49922 430
rect 50038 400 50090 430
rect 50206 400 50258 430
rect 50374 400 50426 430
rect 50542 400 50594 430
rect 50710 400 50762 430
rect 50878 400 50930 430
rect 51046 400 51098 430
rect 51214 400 51266 430
rect 51382 400 51434 430
rect 51550 400 51602 430
rect 51718 400 51770 430
rect 51886 400 51938 430
rect 52054 400 52106 430
rect 52222 400 52274 430
rect 52390 400 52442 430
rect 52558 400 52610 430
rect 52726 400 52778 430
rect 52894 400 52946 430
rect 53062 400 53114 430
rect 53230 400 53282 430
rect 53398 400 53450 430
rect 53566 400 53618 430
rect 53734 400 53786 430
rect 53902 400 53954 430
rect 54070 400 54122 430
rect 54238 400 54290 430
rect 54406 400 54458 430
rect 54574 400 54626 430
rect 54742 400 54794 430
rect 54910 400 54962 430
rect 55078 400 55130 430
rect 55246 400 58842 430
<< obsm3 >>
rect 2233 1554 56135 58422
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
rect 55984 1538 56144 58438
<< labels >>
rlabel metal2 s 1232 59600 1288 60000 6 io_active
port 1 nsew signal input
rlabel metal2 s 1736 59600 1792 60000 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 16856 59600 16912 60000 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 18368 59600 18424 60000 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 19880 59600 19936 60000 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 21392 59600 21448 60000 6 io_in[13]
port 6 nsew signal input
rlabel metal2 s 22904 59600 22960 60000 6 io_in[14]
port 7 nsew signal input
rlabel metal2 s 24416 59600 24472 60000 6 io_in[15]
port 8 nsew signal input
rlabel metal2 s 25928 59600 25984 60000 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 27440 59600 27496 60000 6 io_in[17]
port 10 nsew signal input
rlabel metal2 s 28952 59600 29008 60000 6 io_in[18]
port 11 nsew signal input
rlabel metal2 s 30464 59600 30520 60000 6 io_in[19]
port 12 nsew signal input
rlabel metal2 s 3248 59600 3304 60000 6 io_in[1]
port 13 nsew signal input
rlabel metal2 s 31976 59600 32032 60000 6 io_in[20]
port 14 nsew signal input
rlabel metal2 s 33488 59600 33544 60000 6 io_in[21]
port 15 nsew signal input
rlabel metal2 s 35000 59600 35056 60000 6 io_in[22]
port 16 nsew signal input
rlabel metal2 s 36512 59600 36568 60000 6 io_in[23]
port 17 nsew signal input
rlabel metal2 s 38024 59600 38080 60000 6 io_in[24]
port 18 nsew signal input
rlabel metal2 s 39536 59600 39592 60000 6 io_in[25]
port 19 nsew signal input
rlabel metal2 s 41048 59600 41104 60000 6 io_in[26]
port 20 nsew signal input
rlabel metal2 s 42560 59600 42616 60000 6 io_in[27]
port 21 nsew signal input
rlabel metal2 s 44072 59600 44128 60000 6 io_in[28]
port 22 nsew signal input
rlabel metal2 s 45584 59600 45640 60000 6 io_in[29]
port 23 nsew signal input
rlabel metal2 s 4760 59600 4816 60000 6 io_in[2]
port 24 nsew signal input
rlabel metal2 s 47096 59600 47152 60000 6 io_in[30]
port 25 nsew signal input
rlabel metal2 s 48608 59600 48664 60000 6 io_in[31]
port 26 nsew signal input
rlabel metal2 s 50120 59600 50176 60000 6 io_in[32]
port 27 nsew signal input
rlabel metal2 s 51632 59600 51688 60000 6 io_in[33]
port 28 nsew signal input
rlabel metal2 s 53144 59600 53200 60000 6 io_in[34]
port 29 nsew signal input
rlabel metal2 s 54656 59600 54712 60000 6 io_in[35]
port 30 nsew signal input
rlabel metal2 s 56168 59600 56224 60000 6 io_in[36]
port 31 nsew signal input
rlabel metal2 s 57680 59600 57736 60000 6 io_in[37]
port 32 nsew signal input
rlabel metal2 s 6272 59600 6328 60000 6 io_in[3]
port 33 nsew signal input
rlabel metal2 s 7784 59600 7840 60000 6 io_in[4]
port 34 nsew signal input
rlabel metal2 s 9296 59600 9352 60000 6 io_in[5]
port 35 nsew signal input
rlabel metal2 s 10808 59600 10864 60000 6 io_in[6]
port 36 nsew signal input
rlabel metal2 s 12320 59600 12376 60000 6 io_in[7]
port 37 nsew signal input
rlabel metal2 s 13832 59600 13888 60000 6 io_in[8]
port 38 nsew signal input
rlabel metal2 s 15344 59600 15400 60000 6 io_in[9]
port 39 nsew signal input
rlabel metal2 s 2240 59600 2296 60000 6 io_oeb[0]
port 40 nsew signal output
rlabel metal2 s 17360 59600 17416 60000 6 io_oeb[10]
port 41 nsew signal output
rlabel metal2 s 18872 59600 18928 60000 6 io_oeb[11]
port 42 nsew signal output
rlabel metal2 s 20384 59600 20440 60000 6 io_oeb[12]
port 43 nsew signal output
rlabel metal2 s 21896 59600 21952 60000 6 io_oeb[13]
port 44 nsew signal output
rlabel metal2 s 23408 59600 23464 60000 6 io_oeb[14]
port 45 nsew signal output
rlabel metal2 s 24920 59600 24976 60000 6 io_oeb[15]
port 46 nsew signal output
rlabel metal2 s 26432 59600 26488 60000 6 io_oeb[16]
port 47 nsew signal output
rlabel metal2 s 27944 59600 28000 60000 6 io_oeb[17]
port 48 nsew signal output
rlabel metal2 s 29456 59600 29512 60000 6 io_oeb[18]
port 49 nsew signal output
rlabel metal2 s 30968 59600 31024 60000 6 io_oeb[19]
port 50 nsew signal output
rlabel metal2 s 3752 59600 3808 60000 6 io_oeb[1]
port 51 nsew signal output
rlabel metal2 s 32480 59600 32536 60000 6 io_oeb[20]
port 52 nsew signal output
rlabel metal2 s 33992 59600 34048 60000 6 io_oeb[21]
port 53 nsew signal output
rlabel metal2 s 35504 59600 35560 60000 6 io_oeb[22]
port 54 nsew signal output
rlabel metal2 s 37016 59600 37072 60000 6 io_oeb[23]
port 55 nsew signal output
rlabel metal2 s 38528 59600 38584 60000 6 io_oeb[24]
port 56 nsew signal output
rlabel metal2 s 40040 59600 40096 60000 6 io_oeb[25]
port 57 nsew signal output
rlabel metal2 s 41552 59600 41608 60000 6 io_oeb[26]
port 58 nsew signal output
rlabel metal2 s 43064 59600 43120 60000 6 io_oeb[27]
port 59 nsew signal output
rlabel metal2 s 44576 59600 44632 60000 6 io_oeb[28]
port 60 nsew signal output
rlabel metal2 s 46088 59600 46144 60000 6 io_oeb[29]
port 61 nsew signal output
rlabel metal2 s 5264 59600 5320 60000 6 io_oeb[2]
port 62 nsew signal output
rlabel metal2 s 47600 59600 47656 60000 6 io_oeb[30]
port 63 nsew signal output
rlabel metal2 s 49112 59600 49168 60000 6 io_oeb[31]
port 64 nsew signal output
rlabel metal2 s 50624 59600 50680 60000 6 io_oeb[32]
port 65 nsew signal output
rlabel metal2 s 52136 59600 52192 60000 6 io_oeb[33]
port 66 nsew signal output
rlabel metal2 s 53648 59600 53704 60000 6 io_oeb[34]
port 67 nsew signal output
rlabel metal2 s 55160 59600 55216 60000 6 io_oeb[35]
port 68 nsew signal output
rlabel metal2 s 56672 59600 56728 60000 6 io_oeb[36]
port 69 nsew signal output
rlabel metal2 s 58184 59600 58240 60000 6 io_oeb[37]
port 70 nsew signal output
rlabel metal2 s 6776 59600 6832 60000 6 io_oeb[3]
port 71 nsew signal output
rlabel metal2 s 8288 59600 8344 60000 6 io_oeb[4]
port 72 nsew signal output
rlabel metal2 s 9800 59600 9856 60000 6 io_oeb[5]
port 73 nsew signal output
rlabel metal2 s 11312 59600 11368 60000 6 io_oeb[6]
port 74 nsew signal output
rlabel metal2 s 12824 59600 12880 60000 6 io_oeb[7]
port 75 nsew signal output
rlabel metal2 s 14336 59600 14392 60000 6 io_oeb[8]
port 76 nsew signal output
rlabel metal2 s 15848 59600 15904 60000 6 io_oeb[9]
port 77 nsew signal output
rlabel metal2 s 2744 59600 2800 60000 6 io_out[0]
port 78 nsew signal output
rlabel metal2 s 17864 59600 17920 60000 6 io_out[10]
port 79 nsew signal output
rlabel metal2 s 19376 59600 19432 60000 6 io_out[11]
port 80 nsew signal output
rlabel metal2 s 20888 59600 20944 60000 6 io_out[12]
port 81 nsew signal output
rlabel metal2 s 22400 59600 22456 60000 6 io_out[13]
port 82 nsew signal output
rlabel metal2 s 23912 59600 23968 60000 6 io_out[14]
port 83 nsew signal output
rlabel metal2 s 25424 59600 25480 60000 6 io_out[15]
port 84 nsew signal output
rlabel metal2 s 26936 59600 26992 60000 6 io_out[16]
port 85 nsew signal output
rlabel metal2 s 28448 59600 28504 60000 6 io_out[17]
port 86 nsew signal output
rlabel metal2 s 29960 59600 30016 60000 6 io_out[18]
port 87 nsew signal output
rlabel metal2 s 31472 59600 31528 60000 6 io_out[19]
port 88 nsew signal output
rlabel metal2 s 4256 59600 4312 60000 6 io_out[1]
port 89 nsew signal output
rlabel metal2 s 32984 59600 33040 60000 6 io_out[20]
port 90 nsew signal output
rlabel metal2 s 34496 59600 34552 60000 6 io_out[21]
port 91 nsew signal output
rlabel metal2 s 36008 59600 36064 60000 6 io_out[22]
port 92 nsew signal output
rlabel metal2 s 37520 59600 37576 60000 6 io_out[23]
port 93 nsew signal output
rlabel metal2 s 39032 59600 39088 60000 6 io_out[24]
port 94 nsew signal output
rlabel metal2 s 40544 59600 40600 60000 6 io_out[25]
port 95 nsew signal output
rlabel metal2 s 42056 59600 42112 60000 6 io_out[26]
port 96 nsew signal output
rlabel metal2 s 43568 59600 43624 60000 6 io_out[27]
port 97 nsew signal output
rlabel metal2 s 45080 59600 45136 60000 6 io_out[28]
port 98 nsew signal output
rlabel metal2 s 46592 59600 46648 60000 6 io_out[29]
port 99 nsew signal output
rlabel metal2 s 5768 59600 5824 60000 6 io_out[2]
port 100 nsew signal output
rlabel metal2 s 48104 59600 48160 60000 6 io_out[30]
port 101 nsew signal output
rlabel metal2 s 49616 59600 49672 60000 6 io_out[31]
port 102 nsew signal output
rlabel metal2 s 51128 59600 51184 60000 6 io_out[32]
port 103 nsew signal output
rlabel metal2 s 52640 59600 52696 60000 6 io_out[33]
port 104 nsew signal output
rlabel metal2 s 54152 59600 54208 60000 6 io_out[34]
port 105 nsew signal output
rlabel metal2 s 55664 59600 55720 60000 6 io_out[35]
port 106 nsew signal output
rlabel metal2 s 57176 59600 57232 60000 6 io_out[36]
port 107 nsew signal output
rlabel metal2 s 58688 59600 58744 60000 6 io_out[37]
port 108 nsew signal output
rlabel metal2 s 7280 59600 7336 60000 6 io_out[3]
port 109 nsew signal output
rlabel metal2 s 8792 59600 8848 60000 6 io_out[4]
port 110 nsew signal output
rlabel metal2 s 10304 59600 10360 60000 6 io_out[5]
port 111 nsew signal output
rlabel metal2 s 11816 59600 11872 60000 6 io_out[6]
port 112 nsew signal output
rlabel metal2 s 13328 59600 13384 60000 6 io_out[7]
port 113 nsew signal output
rlabel metal2 s 14840 59600 14896 60000 6 io_out[8]
port 114 nsew signal output
rlabel metal2 s 16352 59600 16408 60000 6 io_out[9]
port 115 nsew signal output
rlabel metal2 s 54824 0 54880 400 6 irq[0]
port 116 nsew signal output
rlabel metal2 s 54992 0 55048 400 6 irq[1]
port 117 nsew signal output
rlabel metal2 s 55160 0 55216 400 6 irq[2]
port 118 nsew signal output
rlabel metal2 s 22568 0 22624 400 6 la_data_in[0]
port 119 nsew signal input
rlabel metal2 s 27608 0 27664 400 6 la_data_in[10]
port 120 nsew signal input
rlabel metal2 s 28112 0 28168 400 6 la_data_in[11]
port 121 nsew signal input
rlabel metal2 s 28616 0 28672 400 6 la_data_in[12]
port 122 nsew signal input
rlabel metal2 s 29120 0 29176 400 6 la_data_in[13]
port 123 nsew signal input
rlabel metal2 s 29624 0 29680 400 6 la_data_in[14]
port 124 nsew signal input
rlabel metal2 s 30128 0 30184 400 6 la_data_in[15]
port 125 nsew signal input
rlabel metal2 s 30632 0 30688 400 6 la_data_in[16]
port 126 nsew signal input
rlabel metal2 s 31136 0 31192 400 6 la_data_in[17]
port 127 nsew signal input
rlabel metal2 s 31640 0 31696 400 6 la_data_in[18]
port 128 nsew signal input
rlabel metal2 s 32144 0 32200 400 6 la_data_in[19]
port 129 nsew signal input
rlabel metal2 s 23072 0 23128 400 6 la_data_in[1]
port 130 nsew signal input
rlabel metal2 s 32648 0 32704 400 6 la_data_in[20]
port 131 nsew signal input
rlabel metal2 s 33152 0 33208 400 6 la_data_in[21]
port 132 nsew signal input
rlabel metal2 s 33656 0 33712 400 6 la_data_in[22]
port 133 nsew signal input
rlabel metal2 s 34160 0 34216 400 6 la_data_in[23]
port 134 nsew signal input
rlabel metal2 s 34664 0 34720 400 6 la_data_in[24]
port 135 nsew signal input
rlabel metal2 s 35168 0 35224 400 6 la_data_in[25]
port 136 nsew signal input
rlabel metal2 s 35672 0 35728 400 6 la_data_in[26]
port 137 nsew signal input
rlabel metal2 s 36176 0 36232 400 6 la_data_in[27]
port 138 nsew signal input
rlabel metal2 s 36680 0 36736 400 6 la_data_in[28]
port 139 nsew signal input
rlabel metal2 s 37184 0 37240 400 6 la_data_in[29]
port 140 nsew signal input
rlabel metal2 s 23576 0 23632 400 6 la_data_in[2]
port 141 nsew signal input
rlabel metal2 s 37688 0 37744 400 6 la_data_in[30]
port 142 nsew signal input
rlabel metal2 s 38192 0 38248 400 6 la_data_in[31]
port 143 nsew signal input
rlabel metal2 s 38696 0 38752 400 6 la_data_in[32]
port 144 nsew signal input
rlabel metal2 s 39200 0 39256 400 6 la_data_in[33]
port 145 nsew signal input
rlabel metal2 s 39704 0 39760 400 6 la_data_in[34]
port 146 nsew signal input
rlabel metal2 s 40208 0 40264 400 6 la_data_in[35]
port 147 nsew signal input
rlabel metal2 s 40712 0 40768 400 6 la_data_in[36]
port 148 nsew signal input
rlabel metal2 s 41216 0 41272 400 6 la_data_in[37]
port 149 nsew signal input
rlabel metal2 s 41720 0 41776 400 6 la_data_in[38]
port 150 nsew signal input
rlabel metal2 s 42224 0 42280 400 6 la_data_in[39]
port 151 nsew signal input
rlabel metal2 s 24080 0 24136 400 6 la_data_in[3]
port 152 nsew signal input
rlabel metal2 s 42728 0 42784 400 6 la_data_in[40]
port 153 nsew signal input
rlabel metal2 s 43232 0 43288 400 6 la_data_in[41]
port 154 nsew signal input
rlabel metal2 s 43736 0 43792 400 6 la_data_in[42]
port 155 nsew signal input
rlabel metal2 s 44240 0 44296 400 6 la_data_in[43]
port 156 nsew signal input
rlabel metal2 s 44744 0 44800 400 6 la_data_in[44]
port 157 nsew signal input
rlabel metal2 s 45248 0 45304 400 6 la_data_in[45]
port 158 nsew signal input
rlabel metal2 s 45752 0 45808 400 6 la_data_in[46]
port 159 nsew signal input
rlabel metal2 s 46256 0 46312 400 6 la_data_in[47]
port 160 nsew signal input
rlabel metal2 s 46760 0 46816 400 6 la_data_in[48]
port 161 nsew signal input
rlabel metal2 s 47264 0 47320 400 6 la_data_in[49]
port 162 nsew signal input
rlabel metal2 s 24584 0 24640 400 6 la_data_in[4]
port 163 nsew signal input
rlabel metal2 s 47768 0 47824 400 6 la_data_in[50]
port 164 nsew signal input
rlabel metal2 s 48272 0 48328 400 6 la_data_in[51]
port 165 nsew signal input
rlabel metal2 s 48776 0 48832 400 6 la_data_in[52]
port 166 nsew signal input
rlabel metal2 s 49280 0 49336 400 6 la_data_in[53]
port 167 nsew signal input
rlabel metal2 s 49784 0 49840 400 6 la_data_in[54]
port 168 nsew signal input
rlabel metal2 s 50288 0 50344 400 6 la_data_in[55]
port 169 nsew signal input
rlabel metal2 s 50792 0 50848 400 6 la_data_in[56]
port 170 nsew signal input
rlabel metal2 s 51296 0 51352 400 6 la_data_in[57]
port 171 nsew signal input
rlabel metal2 s 51800 0 51856 400 6 la_data_in[58]
port 172 nsew signal input
rlabel metal2 s 52304 0 52360 400 6 la_data_in[59]
port 173 nsew signal input
rlabel metal2 s 25088 0 25144 400 6 la_data_in[5]
port 174 nsew signal input
rlabel metal2 s 52808 0 52864 400 6 la_data_in[60]
port 175 nsew signal input
rlabel metal2 s 53312 0 53368 400 6 la_data_in[61]
port 176 nsew signal input
rlabel metal2 s 53816 0 53872 400 6 la_data_in[62]
port 177 nsew signal input
rlabel metal2 s 54320 0 54376 400 6 la_data_in[63]
port 178 nsew signal input
rlabel metal2 s 25592 0 25648 400 6 la_data_in[6]
port 179 nsew signal input
rlabel metal2 s 26096 0 26152 400 6 la_data_in[7]
port 180 nsew signal input
rlabel metal2 s 26600 0 26656 400 6 la_data_in[8]
port 181 nsew signal input
rlabel metal2 s 27104 0 27160 400 6 la_data_in[9]
port 182 nsew signal input
rlabel metal2 s 22736 0 22792 400 6 la_data_out[0]
port 183 nsew signal output
rlabel metal2 s 27776 0 27832 400 6 la_data_out[10]
port 184 nsew signal output
rlabel metal2 s 28280 0 28336 400 6 la_data_out[11]
port 185 nsew signal output
rlabel metal2 s 28784 0 28840 400 6 la_data_out[12]
port 186 nsew signal output
rlabel metal2 s 29288 0 29344 400 6 la_data_out[13]
port 187 nsew signal output
rlabel metal2 s 29792 0 29848 400 6 la_data_out[14]
port 188 nsew signal output
rlabel metal2 s 30296 0 30352 400 6 la_data_out[15]
port 189 nsew signal output
rlabel metal2 s 30800 0 30856 400 6 la_data_out[16]
port 190 nsew signal output
rlabel metal2 s 31304 0 31360 400 6 la_data_out[17]
port 191 nsew signal output
rlabel metal2 s 31808 0 31864 400 6 la_data_out[18]
port 192 nsew signal output
rlabel metal2 s 32312 0 32368 400 6 la_data_out[19]
port 193 nsew signal output
rlabel metal2 s 23240 0 23296 400 6 la_data_out[1]
port 194 nsew signal output
rlabel metal2 s 32816 0 32872 400 6 la_data_out[20]
port 195 nsew signal output
rlabel metal2 s 33320 0 33376 400 6 la_data_out[21]
port 196 nsew signal output
rlabel metal2 s 33824 0 33880 400 6 la_data_out[22]
port 197 nsew signal output
rlabel metal2 s 34328 0 34384 400 6 la_data_out[23]
port 198 nsew signal output
rlabel metal2 s 34832 0 34888 400 6 la_data_out[24]
port 199 nsew signal output
rlabel metal2 s 35336 0 35392 400 6 la_data_out[25]
port 200 nsew signal output
rlabel metal2 s 35840 0 35896 400 6 la_data_out[26]
port 201 nsew signal output
rlabel metal2 s 36344 0 36400 400 6 la_data_out[27]
port 202 nsew signal output
rlabel metal2 s 36848 0 36904 400 6 la_data_out[28]
port 203 nsew signal output
rlabel metal2 s 37352 0 37408 400 6 la_data_out[29]
port 204 nsew signal output
rlabel metal2 s 23744 0 23800 400 6 la_data_out[2]
port 205 nsew signal output
rlabel metal2 s 37856 0 37912 400 6 la_data_out[30]
port 206 nsew signal output
rlabel metal2 s 38360 0 38416 400 6 la_data_out[31]
port 207 nsew signal output
rlabel metal2 s 38864 0 38920 400 6 la_data_out[32]
port 208 nsew signal output
rlabel metal2 s 39368 0 39424 400 6 la_data_out[33]
port 209 nsew signal output
rlabel metal2 s 39872 0 39928 400 6 la_data_out[34]
port 210 nsew signal output
rlabel metal2 s 40376 0 40432 400 6 la_data_out[35]
port 211 nsew signal output
rlabel metal2 s 40880 0 40936 400 6 la_data_out[36]
port 212 nsew signal output
rlabel metal2 s 41384 0 41440 400 6 la_data_out[37]
port 213 nsew signal output
rlabel metal2 s 41888 0 41944 400 6 la_data_out[38]
port 214 nsew signal output
rlabel metal2 s 42392 0 42448 400 6 la_data_out[39]
port 215 nsew signal output
rlabel metal2 s 24248 0 24304 400 6 la_data_out[3]
port 216 nsew signal output
rlabel metal2 s 42896 0 42952 400 6 la_data_out[40]
port 217 nsew signal output
rlabel metal2 s 43400 0 43456 400 6 la_data_out[41]
port 218 nsew signal output
rlabel metal2 s 43904 0 43960 400 6 la_data_out[42]
port 219 nsew signal output
rlabel metal2 s 44408 0 44464 400 6 la_data_out[43]
port 220 nsew signal output
rlabel metal2 s 44912 0 44968 400 6 la_data_out[44]
port 221 nsew signal output
rlabel metal2 s 45416 0 45472 400 6 la_data_out[45]
port 222 nsew signal output
rlabel metal2 s 45920 0 45976 400 6 la_data_out[46]
port 223 nsew signal output
rlabel metal2 s 46424 0 46480 400 6 la_data_out[47]
port 224 nsew signal output
rlabel metal2 s 46928 0 46984 400 6 la_data_out[48]
port 225 nsew signal output
rlabel metal2 s 47432 0 47488 400 6 la_data_out[49]
port 226 nsew signal output
rlabel metal2 s 24752 0 24808 400 6 la_data_out[4]
port 227 nsew signal output
rlabel metal2 s 47936 0 47992 400 6 la_data_out[50]
port 228 nsew signal output
rlabel metal2 s 48440 0 48496 400 6 la_data_out[51]
port 229 nsew signal output
rlabel metal2 s 48944 0 49000 400 6 la_data_out[52]
port 230 nsew signal output
rlabel metal2 s 49448 0 49504 400 6 la_data_out[53]
port 231 nsew signal output
rlabel metal2 s 49952 0 50008 400 6 la_data_out[54]
port 232 nsew signal output
rlabel metal2 s 50456 0 50512 400 6 la_data_out[55]
port 233 nsew signal output
rlabel metal2 s 50960 0 51016 400 6 la_data_out[56]
port 234 nsew signal output
rlabel metal2 s 51464 0 51520 400 6 la_data_out[57]
port 235 nsew signal output
rlabel metal2 s 51968 0 52024 400 6 la_data_out[58]
port 236 nsew signal output
rlabel metal2 s 52472 0 52528 400 6 la_data_out[59]
port 237 nsew signal output
rlabel metal2 s 25256 0 25312 400 6 la_data_out[5]
port 238 nsew signal output
rlabel metal2 s 52976 0 53032 400 6 la_data_out[60]
port 239 nsew signal output
rlabel metal2 s 53480 0 53536 400 6 la_data_out[61]
port 240 nsew signal output
rlabel metal2 s 53984 0 54040 400 6 la_data_out[62]
port 241 nsew signal output
rlabel metal2 s 54488 0 54544 400 6 la_data_out[63]
port 242 nsew signal output
rlabel metal2 s 25760 0 25816 400 6 la_data_out[6]
port 243 nsew signal output
rlabel metal2 s 26264 0 26320 400 6 la_data_out[7]
port 244 nsew signal output
rlabel metal2 s 26768 0 26824 400 6 la_data_out[8]
port 245 nsew signal output
rlabel metal2 s 27272 0 27328 400 6 la_data_out[9]
port 246 nsew signal output
rlabel metal2 s 22904 0 22960 400 6 la_oenb[0]
port 247 nsew signal input
rlabel metal2 s 27944 0 28000 400 6 la_oenb[10]
port 248 nsew signal input
rlabel metal2 s 28448 0 28504 400 6 la_oenb[11]
port 249 nsew signal input
rlabel metal2 s 28952 0 29008 400 6 la_oenb[12]
port 250 nsew signal input
rlabel metal2 s 29456 0 29512 400 6 la_oenb[13]
port 251 nsew signal input
rlabel metal2 s 29960 0 30016 400 6 la_oenb[14]
port 252 nsew signal input
rlabel metal2 s 30464 0 30520 400 6 la_oenb[15]
port 253 nsew signal input
rlabel metal2 s 30968 0 31024 400 6 la_oenb[16]
port 254 nsew signal input
rlabel metal2 s 31472 0 31528 400 6 la_oenb[17]
port 255 nsew signal input
rlabel metal2 s 31976 0 32032 400 6 la_oenb[18]
port 256 nsew signal input
rlabel metal2 s 32480 0 32536 400 6 la_oenb[19]
port 257 nsew signal input
rlabel metal2 s 23408 0 23464 400 6 la_oenb[1]
port 258 nsew signal input
rlabel metal2 s 32984 0 33040 400 6 la_oenb[20]
port 259 nsew signal input
rlabel metal2 s 33488 0 33544 400 6 la_oenb[21]
port 260 nsew signal input
rlabel metal2 s 33992 0 34048 400 6 la_oenb[22]
port 261 nsew signal input
rlabel metal2 s 34496 0 34552 400 6 la_oenb[23]
port 262 nsew signal input
rlabel metal2 s 35000 0 35056 400 6 la_oenb[24]
port 263 nsew signal input
rlabel metal2 s 35504 0 35560 400 6 la_oenb[25]
port 264 nsew signal input
rlabel metal2 s 36008 0 36064 400 6 la_oenb[26]
port 265 nsew signal input
rlabel metal2 s 36512 0 36568 400 6 la_oenb[27]
port 266 nsew signal input
rlabel metal2 s 37016 0 37072 400 6 la_oenb[28]
port 267 nsew signal input
rlabel metal2 s 37520 0 37576 400 6 la_oenb[29]
port 268 nsew signal input
rlabel metal2 s 23912 0 23968 400 6 la_oenb[2]
port 269 nsew signal input
rlabel metal2 s 38024 0 38080 400 6 la_oenb[30]
port 270 nsew signal input
rlabel metal2 s 38528 0 38584 400 6 la_oenb[31]
port 271 nsew signal input
rlabel metal2 s 39032 0 39088 400 6 la_oenb[32]
port 272 nsew signal input
rlabel metal2 s 39536 0 39592 400 6 la_oenb[33]
port 273 nsew signal input
rlabel metal2 s 40040 0 40096 400 6 la_oenb[34]
port 274 nsew signal input
rlabel metal2 s 40544 0 40600 400 6 la_oenb[35]
port 275 nsew signal input
rlabel metal2 s 41048 0 41104 400 6 la_oenb[36]
port 276 nsew signal input
rlabel metal2 s 41552 0 41608 400 6 la_oenb[37]
port 277 nsew signal input
rlabel metal2 s 42056 0 42112 400 6 la_oenb[38]
port 278 nsew signal input
rlabel metal2 s 42560 0 42616 400 6 la_oenb[39]
port 279 nsew signal input
rlabel metal2 s 24416 0 24472 400 6 la_oenb[3]
port 280 nsew signal input
rlabel metal2 s 43064 0 43120 400 6 la_oenb[40]
port 281 nsew signal input
rlabel metal2 s 43568 0 43624 400 6 la_oenb[41]
port 282 nsew signal input
rlabel metal2 s 44072 0 44128 400 6 la_oenb[42]
port 283 nsew signal input
rlabel metal2 s 44576 0 44632 400 6 la_oenb[43]
port 284 nsew signal input
rlabel metal2 s 45080 0 45136 400 6 la_oenb[44]
port 285 nsew signal input
rlabel metal2 s 45584 0 45640 400 6 la_oenb[45]
port 286 nsew signal input
rlabel metal2 s 46088 0 46144 400 6 la_oenb[46]
port 287 nsew signal input
rlabel metal2 s 46592 0 46648 400 6 la_oenb[47]
port 288 nsew signal input
rlabel metal2 s 47096 0 47152 400 6 la_oenb[48]
port 289 nsew signal input
rlabel metal2 s 47600 0 47656 400 6 la_oenb[49]
port 290 nsew signal input
rlabel metal2 s 24920 0 24976 400 6 la_oenb[4]
port 291 nsew signal input
rlabel metal2 s 48104 0 48160 400 6 la_oenb[50]
port 292 nsew signal input
rlabel metal2 s 48608 0 48664 400 6 la_oenb[51]
port 293 nsew signal input
rlabel metal2 s 49112 0 49168 400 6 la_oenb[52]
port 294 nsew signal input
rlabel metal2 s 49616 0 49672 400 6 la_oenb[53]
port 295 nsew signal input
rlabel metal2 s 50120 0 50176 400 6 la_oenb[54]
port 296 nsew signal input
rlabel metal2 s 50624 0 50680 400 6 la_oenb[55]
port 297 nsew signal input
rlabel metal2 s 51128 0 51184 400 6 la_oenb[56]
port 298 nsew signal input
rlabel metal2 s 51632 0 51688 400 6 la_oenb[57]
port 299 nsew signal input
rlabel metal2 s 52136 0 52192 400 6 la_oenb[58]
port 300 nsew signal input
rlabel metal2 s 52640 0 52696 400 6 la_oenb[59]
port 301 nsew signal input
rlabel metal2 s 25424 0 25480 400 6 la_oenb[5]
port 302 nsew signal input
rlabel metal2 s 53144 0 53200 400 6 la_oenb[60]
port 303 nsew signal input
rlabel metal2 s 53648 0 53704 400 6 la_oenb[61]
port 304 nsew signal input
rlabel metal2 s 54152 0 54208 400 6 la_oenb[62]
port 305 nsew signal input
rlabel metal2 s 54656 0 54712 400 6 la_oenb[63]
port 306 nsew signal input
rlabel metal2 s 25928 0 25984 400 6 la_oenb[6]
port 307 nsew signal input
rlabel metal2 s 26432 0 26488 400 6 la_oenb[7]
port 308 nsew signal input
rlabel metal2 s 26936 0 26992 400 6 la_oenb[8]
port 309 nsew signal input
rlabel metal2 s 27440 0 27496 400 6 la_oenb[9]
port 310 nsew signal input
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vdd
port 311 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58438 6 vss
port 312 nsew ground bidirectional
rlabel metal2 s 4760 0 4816 400 6 wb_clk_i
port 313 nsew signal input
rlabel metal2 s 4928 0 4984 400 6 wb_rst_i
port 314 nsew signal input
rlabel metal2 s 5096 0 5152 400 6 wbs_ack_o
port 315 nsew signal output
rlabel metal2 s 5768 0 5824 400 6 wbs_adr_i[0]
port 316 nsew signal input
rlabel metal2 s 11480 0 11536 400 6 wbs_adr_i[10]
port 317 nsew signal input
rlabel metal2 s 11984 0 12040 400 6 wbs_adr_i[11]
port 318 nsew signal input
rlabel metal2 s 12488 0 12544 400 6 wbs_adr_i[12]
port 319 nsew signal input
rlabel metal2 s 12992 0 13048 400 6 wbs_adr_i[13]
port 320 nsew signal input
rlabel metal2 s 13496 0 13552 400 6 wbs_adr_i[14]
port 321 nsew signal input
rlabel metal2 s 14000 0 14056 400 6 wbs_adr_i[15]
port 322 nsew signal input
rlabel metal2 s 14504 0 14560 400 6 wbs_adr_i[16]
port 323 nsew signal input
rlabel metal2 s 15008 0 15064 400 6 wbs_adr_i[17]
port 324 nsew signal input
rlabel metal2 s 15512 0 15568 400 6 wbs_adr_i[18]
port 325 nsew signal input
rlabel metal2 s 16016 0 16072 400 6 wbs_adr_i[19]
port 326 nsew signal input
rlabel metal2 s 6440 0 6496 400 6 wbs_adr_i[1]
port 327 nsew signal input
rlabel metal2 s 16520 0 16576 400 6 wbs_adr_i[20]
port 328 nsew signal input
rlabel metal2 s 17024 0 17080 400 6 wbs_adr_i[21]
port 329 nsew signal input
rlabel metal2 s 17528 0 17584 400 6 wbs_adr_i[22]
port 330 nsew signal input
rlabel metal2 s 18032 0 18088 400 6 wbs_adr_i[23]
port 331 nsew signal input
rlabel metal2 s 18536 0 18592 400 6 wbs_adr_i[24]
port 332 nsew signal input
rlabel metal2 s 19040 0 19096 400 6 wbs_adr_i[25]
port 333 nsew signal input
rlabel metal2 s 19544 0 19600 400 6 wbs_adr_i[26]
port 334 nsew signal input
rlabel metal2 s 20048 0 20104 400 6 wbs_adr_i[27]
port 335 nsew signal input
rlabel metal2 s 20552 0 20608 400 6 wbs_adr_i[28]
port 336 nsew signal input
rlabel metal2 s 21056 0 21112 400 6 wbs_adr_i[29]
port 337 nsew signal input
rlabel metal2 s 7112 0 7168 400 6 wbs_adr_i[2]
port 338 nsew signal input
rlabel metal2 s 21560 0 21616 400 6 wbs_adr_i[30]
port 339 nsew signal input
rlabel metal2 s 22064 0 22120 400 6 wbs_adr_i[31]
port 340 nsew signal input
rlabel metal2 s 7784 0 7840 400 6 wbs_adr_i[3]
port 341 nsew signal input
rlabel metal2 s 8456 0 8512 400 6 wbs_adr_i[4]
port 342 nsew signal input
rlabel metal2 s 8960 0 9016 400 6 wbs_adr_i[5]
port 343 nsew signal input
rlabel metal2 s 9464 0 9520 400 6 wbs_adr_i[6]
port 344 nsew signal input
rlabel metal2 s 9968 0 10024 400 6 wbs_adr_i[7]
port 345 nsew signal input
rlabel metal2 s 10472 0 10528 400 6 wbs_adr_i[8]
port 346 nsew signal input
rlabel metal2 s 10976 0 11032 400 6 wbs_adr_i[9]
port 347 nsew signal input
rlabel metal2 s 5264 0 5320 400 6 wbs_cyc_i
port 348 nsew signal input
rlabel metal2 s 5936 0 5992 400 6 wbs_dat_i[0]
port 349 nsew signal input
rlabel metal2 s 11648 0 11704 400 6 wbs_dat_i[10]
port 350 nsew signal input
rlabel metal2 s 12152 0 12208 400 6 wbs_dat_i[11]
port 351 nsew signal input
rlabel metal2 s 12656 0 12712 400 6 wbs_dat_i[12]
port 352 nsew signal input
rlabel metal2 s 13160 0 13216 400 6 wbs_dat_i[13]
port 353 nsew signal input
rlabel metal2 s 13664 0 13720 400 6 wbs_dat_i[14]
port 354 nsew signal input
rlabel metal2 s 14168 0 14224 400 6 wbs_dat_i[15]
port 355 nsew signal input
rlabel metal2 s 14672 0 14728 400 6 wbs_dat_i[16]
port 356 nsew signal input
rlabel metal2 s 15176 0 15232 400 6 wbs_dat_i[17]
port 357 nsew signal input
rlabel metal2 s 15680 0 15736 400 6 wbs_dat_i[18]
port 358 nsew signal input
rlabel metal2 s 16184 0 16240 400 6 wbs_dat_i[19]
port 359 nsew signal input
rlabel metal2 s 6608 0 6664 400 6 wbs_dat_i[1]
port 360 nsew signal input
rlabel metal2 s 16688 0 16744 400 6 wbs_dat_i[20]
port 361 nsew signal input
rlabel metal2 s 17192 0 17248 400 6 wbs_dat_i[21]
port 362 nsew signal input
rlabel metal2 s 17696 0 17752 400 6 wbs_dat_i[22]
port 363 nsew signal input
rlabel metal2 s 18200 0 18256 400 6 wbs_dat_i[23]
port 364 nsew signal input
rlabel metal2 s 18704 0 18760 400 6 wbs_dat_i[24]
port 365 nsew signal input
rlabel metal2 s 19208 0 19264 400 6 wbs_dat_i[25]
port 366 nsew signal input
rlabel metal2 s 19712 0 19768 400 6 wbs_dat_i[26]
port 367 nsew signal input
rlabel metal2 s 20216 0 20272 400 6 wbs_dat_i[27]
port 368 nsew signal input
rlabel metal2 s 20720 0 20776 400 6 wbs_dat_i[28]
port 369 nsew signal input
rlabel metal2 s 21224 0 21280 400 6 wbs_dat_i[29]
port 370 nsew signal input
rlabel metal2 s 7280 0 7336 400 6 wbs_dat_i[2]
port 371 nsew signal input
rlabel metal2 s 21728 0 21784 400 6 wbs_dat_i[30]
port 372 nsew signal input
rlabel metal2 s 22232 0 22288 400 6 wbs_dat_i[31]
port 373 nsew signal input
rlabel metal2 s 7952 0 8008 400 6 wbs_dat_i[3]
port 374 nsew signal input
rlabel metal2 s 8624 0 8680 400 6 wbs_dat_i[4]
port 375 nsew signal input
rlabel metal2 s 9128 0 9184 400 6 wbs_dat_i[5]
port 376 nsew signal input
rlabel metal2 s 9632 0 9688 400 6 wbs_dat_i[6]
port 377 nsew signal input
rlabel metal2 s 10136 0 10192 400 6 wbs_dat_i[7]
port 378 nsew signal input
rlabel metal2 s 10640 0 10696 400 6 wbs_dat_i[8]
port 379 nsew signal input
rlabel metal2 s 11144 0 11200 400 6 wbs_dat_i[9]
port 380 nsew signal input
rlabel metal2 s 6104 0 6160 400 6 wbs_dat_o[0]
port 381 nsew signal output
rlabel metal2 s 11816 0 11872 400 6 wbs_dat_o[10]
port 382 nsew signal output
rlabel metal2 s 12320 0 12376 400 6 wbs_dat_o[11]
port 383 nsew signal output
rlabel metal2 s 12824 0 12880 400 6 wbs_dat_o[12]
port 384 nsew signal output
rlabel metal2 s 13328 0 13384 400 6 wbs_dat_o[13]
port 385 nsew signal output
rlabel metal2 s 13832 0 13888 400 6 wbs_dat_o[14]
port 386 nsew signal output
rlabel metal2 s 14336 0 14392 400 6 wbs_dat_o[15]
port 387 nsew signal output
rlabel metal2 s 14840 0 14896 400 6 wbs_dat_o[16]
port 388 nsew signal output
rlabel metal2 s 15344 0 15400 400 6 wbs_dat_o[17]
port 389 nsew signal output
rlabel metal2 s 15848 0 15904 400 6 wbs_dat_o[18]
port 390 nsew signal output
rlabel metal2 s 16352 0 16408 400 6 wbs_dat_o[19]
port 391 nsew signal output
rlabel metal2 s 6776 0 6832 400 6 wbs_dat_o[1]
port 392 nsew signal output
rlabel metal2 s 16856 0 16912 400 6 wbs_dat_o[20]
port 393 nsew signal output
rlabel metal2 s 17360 0 17416 400 6 wbs_dat_o[21]
port 394 nsew signal output
rlabel metal2 s 17864 0 17920 400 6 wbs_dat_o[22]
port 395 nsew signal output
rlabel metal2 s 18368 0 18424 400 6 wbs_dat_o[23]
port 396 nsew signal output
rlabel metal2 s 18872 0 18928 400 6 wbs_dat_o[24]
port 397 nsew signal output
rlabel metal2 s 19376 0 19432 400 6 wbs_dat_o[25]
port 398 nsew signal output
rlabel metal2 s 19880 0 19936 400 6 wbs_dat_o[26]
port 399 nsew signal output
rlabel metal2 s 20384 0 20440 400 6 wbs_dat_o[27]
port 400 nsew signal output
rlabel metal2 s 20888 0 20944 400 6 wbs_dat_o[28]
port 401 nsew signal output
rlabel metal2 s 21392 0 21448 400 6 wbs_dat_o[29]
port 402 nsew signal output
rlabel metal2 s 7448 0 7504 400 6 wbs_dat_o[2]
port 403 nsew signal output
rlabel metal2 s 21896 0 21952 400 6 wbs_dat_o[30]
port 404 nsew signal output
rlabel metal2 s 22400 0 22456 400 6 wbs_dat_o[31]
port 405 nsew signal output
rlabel metal2 s 8120 0 8176 400 6 wbs_dat_o[3]
port 406 nsew signal output
rlabel metal2 s 8792 0 8848 400 6 wbs_dat_o[4]
port 407 nsew signal output
rlabel metal2 s 9296 0 9352 400 6 wbs_dat_o[5]
port 408 nsew signal output
rlabel metal2 s 9800 0 9856 400 6 wbs_dat_o[6]
port 409 nsew signal output
rlabel metal2 s 10304 0 10360 400 6 wbs_dat_o[7]
port 410 nsew signal output
rlabel metal2 s 10808 0 10864 400 6 wbs_dat_o[8]
port 411 nsew signal output
rlabel metal2 s 11312 0 11368 400 6 wbs_dat_o[9]
port 412 nsew signal output
rlabel metal2 s 6272 0 6328 400 6 wbs_sel_i[0]
port 413 nsew signal input
rlabel metal2 s 6944 0 7000 400 6 wbs_sel_i[1]
port 414 nsew signal input
rlabel metal2 s 7616 0 7672 400 6 wbs_sel_i[2]
port 415 nsew signal input
rlabel metal2 s 8288 0 8344 400 6 wbs_sel_i[3]
port 416 nsew signal input
rlabel metal2 s 5432 0 5488 400 6 wbs_stb_i
port 417 nsew signal input
rlabel metal2 s 5600 0 5656 400 6 wbs_we_i
port 418 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1462556
string GDS_FILE /opt/gf_180/openlane/user_proj_example/runs/22_12_05_14_45/results/signoff/macro_decap.magic.gds
string GDS_START 48094
<< end >>

