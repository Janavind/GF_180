// This is the unpowered netlist.
module macro_tap (io_active,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    irq,
    la_data_in,
    la_data_out,
    la_oenb,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input io_active;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [2:0] irq;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire net99;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net100;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net101;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net140;
 wire net141;
 wire net137;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net138;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net139;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net164;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net165;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net166;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net167;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net168;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net66;
 wire net67;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net68;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net69;
 wire net97;
 wire net98;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _119_ (.I(net19),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _120_ (.I(_059_),
    .Z(_060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _121_ (.I(_060_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _122_ (.I(net6),
    .Z(_062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _123_ (.A1(net18),
    .A2(_059_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _124_ (.A1(net8),
    .A2(_062_),
    .A3(net7),
    .B(_063_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _125_ (.A1(net9),
    .A2(_064_),
    .Z(_065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _126_ (.A1(net5),
    .A2(_065_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _127_ (.I(net18),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _128_ (.A1(net6),
    .A2(net7),
    .B1(_067_),
    .B2(net19),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _129_ (.A1(net8),
    .A2(_068_),
    .Z(_069_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _130_ (.A1(net4),
    .A2(_069_),
    .Z(_070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _131_ (.I(net3),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _132_ (.I(net7),
    .Z(_072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _133_ (.A1(_067_),
    .A2(net19),
    .B(net6),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _134_ (.A1(_072_),
    .A2(_073_),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _135_ (.A1(_072_),
    .A2(_073_),
    .Z(_075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _136_ (.I(_062_),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _137_ (.A1(_076_),
    .A2(net2),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _138_ (.A1(net7),
    .A2(_071_),
    .A3(_073_),
    .Z(_078_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _139_ (.A1(_071_),
    .A2(_074_),
    .A3(_075_),
    .B1(_077_),
    .B2(_078_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _140_ (.A1(net4),
    .A2(_069_),
    .Z(_080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _141_ (.A1(net5),
    .A2(_065_),
    .B1(_070_),
    .B2(_079_),
    .C(_080_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _142_ (.A1(net9),
    .A2(_063_),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _143_ (.A1(_064_),
    .A2(_082_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _144_ (.A1(_066_),
    .A2(_081_),
    .A3(_083_),
    .Z(_084_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _145_ (.A1(_066_),
    .A2(_081_),
    .B(_083_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _146_ (.A1(_061_),
    .A2(_084_),
    .A3(_085_),
    .Z(_086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _147_ (.I(net21),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _148_ (.I(_087_),
    .Z(_088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _149_ (.I(_088_),
    .Z(_089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _150_ (.A1(net20),
    .A2(_087_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _151_ (.I(net14),
    .Z(_091_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _152_ (.A1(net16),
    .A2(_091_),
    .A3(net15),
    .Z(_092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _153_ (.A1(_090_),
    .A2(_092_),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _154_ (.A1(net17),
    .A2(_093_),
    .Z(_094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _155_ (.A1(net13),
    .A2(_094_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _156_ (.I(net20),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _157_ (.A1(net14),
    .A2(net15),
    .B1(_096_),
    .B2(net21),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _158_ (.A1(net16),
    .A2(_097_),
    .Z(_098_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _159_ (.A1(net12),
    .A2(_098_),
    .Z(_099_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _160_ (.I(net11),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _161_ (.I(net15),
    .Z(_101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _162_ (.A1(_096_),
    .A2(net21),
    .B(net14),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _163_ (.A1(_101_),
    .A2(_102_),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _164_ (.A1(_101_),
    .A2(_102_),
    .Z(_104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _165_ (.I(_091_),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _166_ (.A1(_105_),
    .A2(net10),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _167_ (.A1(net15),
    .A2(_100_),
    .A3(_102_),
    .Z(_107_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _168_ (.A1(_100_),
    .A2(_103_),
    .A3(_104_),
    .B1(_106_),
    .B2(_107_),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _169_ (.A1(net12),
    .A2(_098_),
    .Z(_109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _170_ (.A1(net13),
    .A2(_094_),
    .B1(_099_),
    .B2(_108_),
    .C(_109_),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _171_ (.A1(net17),
    .A2(_092_),
    .B(_090_),
    .ZN(_111_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _172_ (.I(_111_),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _173_ (.A1(_095_),
    .A2(_110_),
    .A3(_112_),
    .Z(_113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _174_ (.A1(_095_),
    .A2(_110_),
    .B(_112_),
    .ZN(_114_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _175_ (.A1(_089_),
    .A2(_113_),
    .A3(_114_),
    .Z(_115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _176_ (.I(net1),
    .Z(_116_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _177_ (.A1(_089_),
    .A2(_116_),
    .A3(_113_),
    .A4(_114_),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _178_ (.A1(_061_),
    .A2(_116_),
    .A3(_084_),
    .A4(_085_),
    .ZN(_118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _179_ (.A1(_086_),
    .A2(_115_),
    .B1(_117_),
    .B2(_118_),
    .ZN(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _180_ (.I(_117_),
    .ZN(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _181_ (.I(_118_),
    .ZN(net32));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _182_ (.A1(_062_),
    .A2(net2),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _183_ (.A1(_062_),
    .A2(net2),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _184_ (.I(net18),
    .Z(_002_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _185_ (.A1(_002_),
    .A2(_060_),
    .B(_000_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _186_ (.A1(_060_),
    .A2(_000_),
    .B1(_001_),
    .B2(_003_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _187_ (.A1(_091_),
    .A2(net10),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _188_ (.A1(_091_),
    .A2(net10),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _189_ (.I(net20),
    .Z(_007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _190_ (.A1(_007_),
    .A2(_088_),
    .B(_005_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _191_ (.A1(_088_),
    .A2(_005_),
    .B1(_006_),
    .B2(_008_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _192_ (.I(net1),
    .Z(_010_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _193_ (.A1(_010_),
    .A2(_009_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _194_ (.I(_011_),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _195_ (.A1(_010_),
    .A2(_004_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _196_ (.I(_012_),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _197_ (.A1(net23),
    .A2(net27),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _198_ (.A1(_004_),
    .A2(_009_),
    .B(_013_),
    .ZN(net33));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _199_ (.A1(_077_),
    .A2(_078_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _200_ (.A1(_072_),
    .A2(_002_),
    .B(net3),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _201_ (.A1(_072_),
    .A2(_002_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _202_ (.A1(_015_),
    .A2(_016_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _203_ (.I(net19),
    .Z(_018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _204_ (.I0(_014_),
    .I1(_017_),
    .S(_018_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _205_ (.A1(_106_),
    .A2(_107_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _206_ (.A1(_101_),
    .A2(_007_),
    .B(net11),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _207_ (.A1(_101_),
    .A2(_007_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _208_ (.A1(_021_),
    .A2(_022_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _209_ (.I(net21),
    .Z(_024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _210_ (.I0(_020_),
    .I1(_023_),
    .S(_024_),
    .Z(_025_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _211_ (.A1(_010_),
    .A2(_025_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _212_ (.I(_026_),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _213_ (.A1(_010_),
    .A2(_019_),
    .Z(_027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _214_ (.I(_027_),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _215_ (.A1(net24),
    .A2(net28),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _216_ (.A1(_019_),
    .A2(_025_),
    .B(_028_),
    .ZN(net34));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _217_ (.A1(_070_),
    .A2(_079_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _218_ (.I(_002_),
    .Z(_030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _219_ (.A1(_030_),
    .A2(net4),
    .B(_060_),
    .C(net8),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _220_ (.A1(_030_),
    .A2(_061_),
    .A3(net4),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _221_ (.A1(_061_),
    .A2(_029_),
    .B(_031_),
    .C(_032_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _222_ (.A1(_099_),
    .A2(_108_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _223_ (.I(_007_),
    .Z(_035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _224_ (.A1(_035_),
    .A2(net12),
    .B(_088_),
    .C(net16),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _225_ (.A1(_035_),
    .A2(_089_),
    .A3(net12),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _226_ (.A1(_089_),
    .A2(_034_),
    .B(_036_),
    .C(_037_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _227_ (.I(_116_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _228_ (.A1(_033_),
    .A2(_038_),
    .B(_039_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _229_ (.A1(_033_),
    .A2(_038_),
    .B(_040_),
    .ZN(net35));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _230_ (.A1(_070_),
    .A2(_079_),
    .B(_080_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _231_ (.A1(net5),
    .A2(_065_),
    .A3(_041_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _232_ (.A1(net9),
    .A2(_030_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _233_ (.A1(net9),
    .A2(_030_),
    .B(net5),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _234_ (.A1(_043_),
    .A2(_044_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _235_ (.I0(_042_),
    .I1(_045_),
    .S(_018_),
    .Z(_046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _236_ (.A1(_099_),
    .A2(_108_),
    .B(_109_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _237_ (.A1(net13),
    .A2(_094_),
    .A3(_047_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _238_ (.A1(net17),
    .A2(_035_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _239_ (.A1(net17),
    .A2(_035_),
    .B(net13),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _240_ (.A1(_049_),
    .A2(_050_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _241_ (.I0(_048_),
    .I1(_051_),
    .S(_024_),
    .Z(_052_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _242_ (.A1(_024_),
    .A2(_049_),
    .A3(_050_),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _243_ (.A1(_024_),
    .A2(_048_),
    .B(_053_),
    .C(_116_),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _244_ (.A1(_018_),
    .A2(_043_),
    .A3(_044_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _245_ (.A1(_018_),
    .A2(_042_),
    .B(_055_),
    .C(_039_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _246_ (.A1(_046_),
    .A2(_052_),
    .B1(_054_),
    .B2(_056_),
    .ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _247_ (.A1(_039_),
    .A2(_038_),
    .Z(_057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _248_ (.I(_057_),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _249_ (.I(_054_),
    .ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _250_ (.A1(_039_),
    .A2(_033_),
    .Z(_058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _251_ (.I(_058_),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _252_ (.I(_056_),
    .ZN(net30));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_38 (.ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_39 (.ZN(net39));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_40 (.ZN(net40));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_41 (.ZN(net41));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_42 (.ZN(net42));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_43 (.ZN(net43));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_44 (.ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_45 (.ZN(net45));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_46 (.ZN(net46));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_47 (.ZN(net47));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_48 (.ZN(net48));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_49 (.ZN(net49));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_50 (.ZN(net50));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_51 (.ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_52 (.ZN(net52));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_53 (.ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_54 (.ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_89 (.ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_90 (.ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_91 (.ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_93 (.ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_94 (.ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_96 (.ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_97 (.ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_98 (.ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_99 (.ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_100 (.ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_101 (.ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_102 (.ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_103 (.ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_104 (.ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_105 (.ZN(net105));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_106 (.ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_107 (.ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_108 (.ZN(net108));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_109 (.ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_110 (.ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_111 (.ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_112 (.ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_113 (.ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_114 (.ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_115 (.ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_116 (.ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_117 (.ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_118 (.ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_119 (.ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_120 (.ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_121 (.ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_122 (.ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_123 (.ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_124 (.ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_125 (.ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_133 (.ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_134 (.ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_135 (.ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_136 (.ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_137 (.ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_138 (.ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_139 (.ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_140 (.ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_141 (.ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_142 (.ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_143 (.ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_144 (.ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_145 (.ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_146 (.ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_147 (.ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_148 (.ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_149 (.ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_150 (.ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_151 (.ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_152 (.ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_153 (.ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_154 (.ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_155 (.ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_156 (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_161 (.ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_162 (.ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_163 (.ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_164 (.ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_165 (.ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_166 (.ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_167 (.ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_168 (.ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_169 (.ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_170 (.ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_171 (.ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_172 (.ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_173 (.ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_174 (.ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_175 (.ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_176 (.ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_177 (.ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_178 (.ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_179 (.ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_180 (.ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_181 (.ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_182 (.ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_183 (.ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_184 (.ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_185 (.ZN(net185));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_186 (.ZN(net186));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_187 (.ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_188 (.ZN(net188));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_189 (.ZN(net189));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_190 (.ZN(net190));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_191 (.ZN(net191));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_192 (.ZN(net192));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_193 (.ZN(net193));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_194 (.ZN(net194));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_195 (.ZN(net195));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_196 (.ZN(net196));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_197 (.ZN(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__218__I (.I(_002_));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(io_active),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input2 (.I(io_in[18]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(io_in[19]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(io_in[20]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input5 (.I(io_in[21]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input6 (.I(io_in[22]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(io_in[23]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input8 (.I(io_in[24]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input9 (.I(io_in[25]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input10 (.I(io_in[26]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input11 (.I(io_in[27]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(io_in[28]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input13 (.I(io_in[29]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input14 (.I(io_in[30]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input15 (.I(io_in[31]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input16 (.I(io_in[32]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input17 (.I(io_in[33]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input18 (.I(io_in[34]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(io_in[35]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input20 (.I(io_in[36]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input21 (.I(io_in[37]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net29),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output31 (.I(net31),
    .Z(io_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net33),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output36 (.I(net36),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__tiel macro_tap_37 (.ZN(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__201__A2 (.I(_002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__200__A2 (.I(_002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__185__A1 (.I(_002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__198__A1 (.I(_004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__195__A2 (.I(_004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__198__A2 (.I(_009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__193__A2 (.I(_009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__243__A1 (.I(_024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__242__A1 (.I(_024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__241__S (.I(_024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__210__S (.I(_024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__216__A2 (.I(_025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__211__A2 (.I(_025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__233__A2 (.I(_030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__232__A2 (.I(_030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__220__A1 (.I(_030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__219__A1 (.I(_030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__247__A2 (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__229__A2 (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__228__A2 (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__245__A2 (.I(_042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__235__I0 (.I(_042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__246__A2 (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__249__I (.I(_054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__246__B1 (.I(_054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__183__A1 (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__182__A1 (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__136__I (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__124__A2 (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__138__A3 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__135__A2 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__134__A2 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__199__A1 (.I(_077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__139__B1 (.I(_077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__171__B (.I(_090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__153__A1 (.I(_090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__188__A1 (.I(_091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__187__A1 (.I(_091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__165__I (.I(_091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__152__A2 (.I(_091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__243__C (.I(_116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__227__I (.I(_116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__178__A2 (.I(_116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__177__A2 (.I(_116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__180__I (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__179__B1 (.I(_117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__181__I (.I(_118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__179__B2 (.I(_118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_active));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_in[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(io_in[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(io_in[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(io_in[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(io_in[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(io_in[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(io_in[32]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(io_in[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(io_in[34]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(io_in[35]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(io_in[36]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(io_in[37]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__192__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__176__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__183__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__182__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__137__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__233__B (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__231__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__141__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__126__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__138__A1 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__132__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__128__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__124__A3 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__219__C (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__129__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__124__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__233__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__232__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__142__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__125__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__225__A3 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__224__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__169__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__159__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__239__B (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__237__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__170__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__155__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__167__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__161__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__157__A2 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__152__A3 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__224__C (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__158__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__152__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__239__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__238__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__171__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__154__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__184__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__127__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__123__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__203__I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__133__A2 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__128__B2 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__119__I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__189__I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__156__I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__150__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__209__I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__162__A2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__157__B2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__147__I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__215__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_687 ();
 assign io_oeb[0] = net98;
 assign io_oeb[10] = net108;
 assign io_oeb[11] = net109;
 assign io_oeb[12] = net110;
 assign io_oeb[13] = net111;
 assign io_oeb[14] = net112;
 assign io_oeb[15] = net113;
 assign io_oeb[16] = net114;
 assign io_oeb[17] = net115;
 assign io_oeb[18] = net116;
 assign io_oeb[19] = net117;
 assign io_oeb[1] = net99;
 assign io_oeb[20] = net118;
 assign io_oeb[21] = net119;
 assign io_oeb[22] = net120;
 assign io_oeb[23] = net121;
 assign io_oeb[24] = net122;
 assign io_oeb[25] = net123;
 assign io_oeb[26] = net124;
 assign io_oeb[27] = net125;
 assign io_oeb[28] = net126;
 assign io_oeb[29] = net127;
 assign io_oeb[2] = net100;
 assign io_oeb[30] = net128;
 assign io_oeb[31] = net129;
 assign io_oeb[32] = net130;
 assign io_oeb[33] = net131;
 assign io_oeb[34] = net132;
 assign io_oeb[35] = net133;
 assign io_oeb[36] = net134;
 assign io_oeb[37] = net135;
 assign io_oeb[3] = net101;
 assign io_oeb[4] = net102;
 assign io_oeb[5] = net103;
 assign io_oeb[6] = net104;
 assign io_oeb[7] = net105;
 assign io_oeb[8] = net106;
 assign io_oeb[9] = net107;
 assign io_out[18] = net139;
 assign io_out[19] = net140;
 assign io_out[1] = net136;
 assign io_out[20] = net141;
 assign io_out[21] = net142;
 assign io_out[22] = net143;
 assign io_out[23] = net144;
 assign io_out[24] = net145;
 assign io_out[25] = net146;
 assign io_out[26] = net147;
 assign io_out[27] = net148;
 assign io_out[28] = net149;
 assign io_out[29] = net150;
 assign io_out[2] = net137;
 assign io_out[30] = net151;
 assign io_out[31] = net152;
 assign io_out[32] = net153;
 assign io_out[33] = net154;
 assign io_out[34] = net155;
 assign io_out[35] = net156;
 assign io_out[36] = net157;
 assign io_out[37] = net158;
 assign io_out[3] = net138;
 assign irq[0] = net159;
 assign irq[1] = net160;
 assign irq[2] = net161;
 assign la_data_out[0] = net162;
 assign la_data_out[10] = net172;
 assign la_data_out[11] = net173;
 assign la_data_out[12] = net174;
 assign la_data_out[13] = net175;
 assign la_data_out[14] = net176;
 assign la_data_out[15] = net177;
 assign la_data_out[16] = net178;
 assign la_data_out[17] = net179;
 assign la_data_out[18] = net180;
 assign la_data_out[19] = net181;
 assign la_data_out[1] = net163;
 assign la_data_out[20] = net182;
 assign la_data_out[21] = net183;
 assign la_data_out[22] = net184;
 assign la_data_out[23] = net185;
 assign la_data_out[24] = net186;
 assign la_data_out[25] = net187;
 assign la_data_out[26] = net188;
 assign la_data_out[27] = net189;
 assign la_data_out[28] = net190;
 assign la_data_out[29] = net191;
 assign la_data_out[2] = net164;
 assign la_data_out[30] = net192;
 assign la_data_out[31] = net193;
 assign la_data_out[32] = net194;
 assign la_data_out[33] = net195;
 assign la_data_out[34] = net196;
 assign la_data_out[35] = net197;
 assign la_data_out[36] = net37;
 assign la_data_out[37] = net38;
 assign la_data_out[38] = net39;
 assign la_data_out[39] = net40;
 assign la_data_out[3] = net165;
 assign la_data_out[40] = net41;
 assign la_data_out[41] = net42;
 assign la_data_out[42] = net43;
 assign la_data_out[43] = net44;
 assign la_data_out[44] = net45;
 assign la_data_out[45] = net46;
 assign la_data_out[46] = net47;
 assign la_data_out[47] = net48;
 assign la_data_out[48] = net49;
 assign la_data_out[49] = net50;
 assign la_data_out[4] = net166;
 assign la_data_out[50] = net51;
 assign la_data_out[51] = net52;
 assign la_data_out[52] = net53;
 assign la_data_out[53] = net54;
 assign la_data_out[54] = net55;
 assign la_data_out[55] = net56;
 assign la_data_out[56] = net57;
 assign la_data_out[57] = net58;
 assign la_data_out[58] = net59;
 assign la_data_out[59] = net60;
 assign la_data_out[5] = net167;
 assign la_data_out[60] = net61;
 assign la_data_out[61] = net62;
 assign la_data_out[62] = net63;
 assign la_data_out[63] = net64;
 assign la_data_out[6] = net168;
 assign la_data_out[7] = net169;
 assign la_data_out[8] = net170;
 assign la_data_out[9] = net171;
 assign wbs_ack_o = net65;
 assign wbs_dat_o[0] = net66;
 assign wbs_dat_o[10] = net76;
 assign wbs_dat_o[11] = net77;
 assign wbs_dat_o[12] = net78;
 assign wbs_dat_o[13] = net79;
 assign wbs_dat_o[14] = net80;
 assign wbs_dat_o[15] = net81;
 assign wbs_dat_o[16] = net82;
 assign wbs_dat_o[17] = net83;
 assign wbs_dat_o[18] = net84;
 assign wbs_dat_o[19] = net85;
 assign wbs_dat_o[1] = net67;
 assign wbs_dat_o[20] = net86;
 assign wbs_dat_o[21] = net87;
 assign wbs_dat_o[22] = net88;
 assign wbs_dat_o[23] = net89;
 assign wbs_dat_o[24] = net90;
 assign wbs_dat_o[25] = net91;
 assign wbs_dat_o[26] = net92;
 assign wbs_dat_o[27] = net93;
 assign wbs_dat_o[28] = net94;
 assign wbs_dat_o[29] = net95;
 assign wbs_dat_o[2] = net68;
 assign wbs_dat_o[30] = net96;
 assign wbs_dat_o[31] = net97;
 assign wbs_dat_o[3] = net69;
 assign wbs_dat_o[4] = net70;
 assign wbs_dat_o[5] = net71;
 assign wbs_dat_o[6] = net72;
 assign wbs_dat_o[7] = net73;
 assign wbs_dat_o[8] = net74;
 assign wbs_dat_o[9] = net75;
endmodule

