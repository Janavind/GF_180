* NGSPICE file created from macro_decap8.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

.subckt macro_decap8 io_active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ irq[0] irq[1] irq[2] la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12]
+ la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18]
+ la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23]
+ la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29]
+ la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34]
+ la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3]
+ la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45]
+ la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50]
+ la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56]
+ la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61]
+ la_data_in[62] la_data_in[63] la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9]
+ la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6]
+ la_data_out[7] la_data_out[8] la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18]
+ la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24]
+ la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30]
+ la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37]
+ la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43]
+ la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4]
+ la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56]
+ la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62]
+ la_oenb[63] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] vdd vss wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_85_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XANTENNA__249__I _054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_93_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_87_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_200_ _072_ _002_ net3 _015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_83_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_131_ net3 _071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_74_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_16
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XANTENNA__162__A2 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_56_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xmacro_decap8_125 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_147 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_158 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_103 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_136 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_114 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_65_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_38_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmacro_decap8_169 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_53_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__135__A2 _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_29_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_89_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput31 net31 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_86_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_93_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_58_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__180__I _117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_70_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_77_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__238__A1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_52_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XANTENNA__229__A1 _033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_130_ net4 _069_ _070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_84_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_65_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmacro_decap8_137 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_104 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_148 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_126 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_115 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_159 irq[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_79_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_50_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input11_I io_in[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xoutput32 net32 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input3_I io_in[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_85_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_85_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_91_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_9_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__247__A2 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XANTENNA__183__A1 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__229__A2 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_189_ net20 _007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__138__A1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_93_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_93_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XANTENNA__129__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmacro_decap8_105 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_116 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xmacro_decap8_138 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_127 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_149 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XANTENNA__233__B net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
Xoutput33 net33 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput22 net22 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_50_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_31_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_89_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XANTENNA__189__I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_91_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_9_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_92_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_188_ _091_ net10 _006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_65_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_47_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xmacro_decap8_106 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_128 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_139 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_117 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_71_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput23 net23 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput34 net34 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_88_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_82_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_85_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_64_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_46_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__239__B net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_77_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_51_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_93_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_187_ _091_ net10 _005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_87_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__138__A3 _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_86_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_62_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_239_ net17 _035_ net13 _050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xmacro_decap8_129 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_107 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_118 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_92_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput24 net24 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput35 net35 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_88_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__201__A2 _002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_85_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_91_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_9_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input1_I io_active vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_82_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__210__S _024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_92_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__159__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_83_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_186_ _060_ _000_ _001_ _003_ _004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_65_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_238_ net17 _035_ _049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_169_ net12 _098_ _109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_92_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmacro_decap8_108 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_119 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_80_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_61_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmacro_decap8_90 wbs_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_43_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_89_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput25 net25 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput36 net36 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_88_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_25_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XANTENNA__195__A2 _004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_89_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_13_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__177__A2 _116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_92_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_60_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_87_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output33_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_185_ _002_ _060_ _000_ _003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XANTENNA__231__A1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_168_ _100_ _103_ _104_ _106_ _107_ _108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_237_ net13 _094_ _047_ _048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmacro_decap8_109 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xmacro_decap8_80 wbs_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_91 wbs_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_88_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_80_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput26 net26 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_88_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_31_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XANTENNA__203__I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_81_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_89_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_13_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_63_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_45_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_87_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_184_ net18 _002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_2_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_16
XFILLER_92_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_60_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_86_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_236_ _099_ _108_ _109_ _047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_167_ net15 _100_ _102_ _107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_92_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
Xmacro_decap8_70 wbs_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_81 wbs_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_92 wbs_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_88_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_219_ _030_ net4 _060_ net8 _031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_93_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xoutput27 net27 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_88_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__198__A1 _004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_1_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_77_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XANTENNA__209__I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_252_ _056_ net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__119__I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_183_ _062_ net2 _001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_1_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_92_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_93_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_86_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_55_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_235_ _042_ _045_ _018_ _046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_70_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_166_ _105_ net10 _106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_61_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
Xmacro_decap8_60 la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_71 wbs_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_82 wbs_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_93 wbs_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_88_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XANTENNA_input18_I io_in[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_37_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_52_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__132__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_149_ _088_ _089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_218_ _002_ _030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_19_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_61_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_34_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput28 net28 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__198__A2 _009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_25_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__127__I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_90_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_16
XFILLER_90_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_31_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_72_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_13_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_54_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_86_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_86_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XANTENNA__243__A1 _024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_182_ _062_ net2 _000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_251_ _058_ net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_77_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output31_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_165_ _091_ _105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_234_ _043_ _044_ _045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_92_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmacro_decap8_61 la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_50 la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_72 wbs_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_83 wbs_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_94 wbs_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_148_ _087_ _088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_217_ _070_ _079_ _029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xoutput29 net29 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_25_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_90_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_85_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_39_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_89_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_5_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_86_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_54_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_250_ _039_ _033_ _058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_181_ _118_ net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__170__A1 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_86_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output24_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__216__A2 _025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_233_ net9 _030_ net5 _044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_164_ _101_ _102_ _104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__152__A1 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
Xmacro_decap8_62 la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_51 la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_40 la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_73 wbs_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_84 wbs_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_95 wbs_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_88_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_87_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_147_ net21 _087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_216_ _019_ _025_ _028_ net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__125__A1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_85_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_89_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_75_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__246__B1 _054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_5_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_180_ _117_ net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_92_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_73_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XANTENNA__225__A3 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_232_ net9 _030_ _043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_163_ _101_ _102_ _103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_73_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmacro_decap8_63 la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_52 la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_41 la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_96 wbs_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_74 wbs_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_85 wbs_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__134__A2 _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_215_ net24 net28 _028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_146_ _061_ _084_ _085_ _086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_19_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input16_I io_in[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_129_ net8 _068_ _069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input8_I io_in[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_16
XFILLER_90_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_60_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XANTENNA__237__A1 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XANTENNA__228__A1 _033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_86_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_89_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_162_ _096_ net21 net14 _102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_231_ net5 _065_ _041_ _042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XANTENNA__152__A3 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmacro_decap8_64 la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_53 la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_42 la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_97 wbs_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_75 wbs_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_86 wbs_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xinput1 io_active net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_83_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_91_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_214_ _027_ net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_145_ _066_ _081_ _083_ _085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_93_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_19_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_40_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_128_ net6 net7 _067_ net19 _068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_93_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_84_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_84_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__246__A2 _052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XANTENNA__181__I _118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__182__A1 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_86_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__228__A2 _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_89_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__176__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XANTENNA__155__A1 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_161_ net15 _101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_230_ _070_ _079_ _080_ _041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_61_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmacro_decap8_43 la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_98 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__128__B2 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmacro_decap8_54 la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_65 wbs_ack_o vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_76 wbs_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_87 wbs_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
Xinput2 io_in[18] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output22_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_213_ _010_ _019_ _027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_144_ _066_ _081_ _083_ _084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_88_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_87_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__184__I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_127_ net18 _067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input21_I io_in[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_21_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_85_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_16
XFILLER_76_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_1_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_73_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__192__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_55_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_160_ net11 _100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
Xmacro_decap8_55 la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_44 la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_66 wbs_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmacro_decap8_99 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__128__A2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmacro_decap8_77 wbs_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_88 wbs_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xinput3 io_in[19] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_91_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_37_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_87_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_87_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_212_ _026_ net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_143_ _064_ _082_ _083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_126_ net5 _065_ _066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input14_I io_in[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_16
XFILLER_72_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_79_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I io_in[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_89_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_91_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XTAP_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_85_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_41_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_70_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_92_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xmacro_decap8_56 la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_45 la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_67 wbs_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_78 wbs_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_89 wbs_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 io_in[20] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_52_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_211_ _010_ _025_ _026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_142_ net9 _063_ _082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_92_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_87_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_90_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_125_ net9 _064_ _065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__200__A2 _002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__185__A1 _002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_72_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__167__A1 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_91_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__158__A1 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_1_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_16
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
Xmacro_decap8_57 la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_46 la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_68 wbs_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_79 wbs_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xinput5 io_in[21] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_210_ _020_ _023_ _024_ _025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_141_ net5 _065_ _070_ _079_ _080_ _081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_70_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_51_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_93_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_92_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_33_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_124_ net8 _062_ net7 _063_ _064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_93_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_15_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_21_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_90_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_12_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_79_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_85_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XANTENNA__171__B _090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_67_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_89_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_85_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xmacro_decap8_58 la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_47 la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_69 wbs_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
Xinput6 io_in[22] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_91_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_87_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_140_ net4 _069_ _080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_93_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_84_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_87_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_123_ net18 _059_ _063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_66_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
Xinput20 io_in[36] net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_84_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__179__B1 _117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_21_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_71_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input12_I io_in[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_91_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input4_I io_in[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_64_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
Xmacro_decap8_48 la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_37 la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_59 la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xinput7 io_in[23] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_199_ _077_ _078_ _014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__197__A1 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_122_ net6 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xinput10 io_in[26] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput21 io_in[37] net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_84_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XANTENNA__179__B2 _118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_81_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_1_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_91_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_82_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_63_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
Xmacro_decap8_49 la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_38 la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xinput8 io_in[24] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_1_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_45_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_60_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_92_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_27_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_198_ _004_ _009_ _013_ net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_92_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_121_ _060_ _061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_15_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput11 io_in[27] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_80_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_21_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_62_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XANTENNA__241__S _024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_81_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_85_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XANTENNA__242__A1 _024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__233__A1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XANTENNA__215__A1 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmacro_decap8_39 la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xinput9 io_in[25] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_51_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_92_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_197_ net23 net27 _013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_120_ _059_ _060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_93_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_15_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput12 io_in[28] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_249_ _054_ net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_84_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XANTENNA__218__I _002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_7_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_89_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XANTENNA_input10_I io_in[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_88_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XANTENNA__224__A2 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input2_I io_in[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XANTENNA__136__I _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__142__A1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_87_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_196_ _012_ net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__124__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_92_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_93_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput13 io_in[29] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_179_ _086_ _115_ _117_ _118_ net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_248_ _057_ net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_88_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_79_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_90_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_81_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_57_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_72_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_90_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_54_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_1_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_36_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__133__A2 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output34_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__147__I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_27_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_195_ _010_ _004_ _012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__124__A2 _062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_33_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
Xinput14 io_in[30] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_247_ _039_ _038_ _057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_15_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_178_ _061_ _116_ _084_ _085_ _118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_56_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_93_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_92_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_38_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_88_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_79_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_50_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_1_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_16
XFILLER_0_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_90_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_91_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_27_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_194_ _011_ net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__124__A3 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_77_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xinput15 io_in[31] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_246_ _046_ _052_ _054_ _056_ net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_177_ _089_ _116_ _113_ _114_ _117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_92_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_88_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_74_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_229_ _033_ _038_ _040_ net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_7_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_93_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_88_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_88_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_85_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_88_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_16
XFILLER_0_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__154__A1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_89_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_16
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
Xmacro_decap8_190 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_51_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_193_ _010_ _009_ _011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
Xinput16 io_in[32] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_245_ _018_ _042_ _055_ _039_ _056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_176_ net1 _116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_92_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input19_I io_in[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_93_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_228_ _033_ _038_ _039_ _040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_159_ net12 _098_ _099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_7_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_93_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_90_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_48_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_63_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_16
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_16
XFILLER_91_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_45_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmacro_decap8_191 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_180 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_86_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_27_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_192_ net1 _010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_89_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_87_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output32_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_244_ _018_ _043_ _044_ _055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xinput17 io_in[33] net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_175_ _089_ _113_ _114_ _115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_93_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_62_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_227_ _116_ _039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_158_ net16 _097_ _098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__239__A1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_93_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_44_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_88_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_90_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmacro_decap8_170 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_60_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmacro_decap8_192 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_181 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_191_ _088_ _005_ _006_ _008_ _009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_1_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_16
XFILLER_92_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_86_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput18 io_in[34] net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_243_ _024_ _048_ _053_ _116_ _054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_174_ _095_ _110_ _112_ _114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_92_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_68_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__224__C net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_157_ net14 net15 _096_ net21 _097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_226_ _089_ _034_ _036_ _037_ _038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_7_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__219__C net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_209_ net21 _024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__157__B2 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_93_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_63_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
Xmacro_decap8_160 irq[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_193 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_182 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_171 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_86_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_190_ _007_ _088_ _005_ _008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_89_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_41_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xinput19 io_in[35] net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_242_ _024_ _049_ _050_ _053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_173_ _095_ _110_ _112_ _113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_23_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_93_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_92_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XANTENNA__193__A2 _009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_87_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_156_ net20 _096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_225_ _035_ _089_ net12 _037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_11_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XANTENNA_input17_I io_in[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_75_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__157__A2 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_208_ _021_ _022_ _023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_139_ _071_ _074_ _075_ _077_ _078_ _079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_85_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input9_I io_in[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_57_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_40_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_81_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmacro_decap8_150 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmacro_decap8_161 irq[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_194 la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_183 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_172 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_63_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_90_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_89_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__243__C _116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_241_ _048_ _051_ _024_ _052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_172_ _111_ _112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_56_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_87_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_224_ _035_ net12 _088_ net16 _036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
X_155_ net13 _094_ _095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_11_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_61_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_88_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_207_ _101_ _007_ _022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_138_ net7 _071_ _073_ _078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_1_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_72_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_79_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_90_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_54_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_89_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_89_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmacro_decap8_151 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_140 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xmacro_decap8_195 la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_184 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_173 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_162 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__211__A2 _025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_89_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_92_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_240_ _049_ _050_ _051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_171_ net17 _092_ _090_ _111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_93_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_92_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XANTENNA_output23_I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_223_ _007_ _035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__169__A1 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_154_ net17 _093_ _094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_88_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_75_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_137_ _076_ net2 _077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_206_ _101_ _007_ net11 _021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_84_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_89_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xmacro_decap8_130 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_152 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_141 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_72_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_53_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
Xmacro_decap8_196 la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_185 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_174 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_163 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_35_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_16
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_17_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_32_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_170_ net13 _094_ _099_ _108_ _109_ _110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_23_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XANTENNA__178__A2 _116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_153_ _090_ _092_ _093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_222_ _099_ _108_ _034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_11_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_93_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_92_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_52_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_87_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_205_ _106_ _107_ _020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_136_ _062_ _076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XANTENNA_input15_I io_in[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__232__A1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_119_ net19 _059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input7_I io_in[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_16
Xmacro_decap8_131 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_153 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_120 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_142 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmacro_decap8_186 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_175 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_164 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xmacro_decap8_197 la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_90_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_16
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_41_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_23_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_55_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_152_ net16 _091_ net15 _092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_221_ _061_ _029_ _031_ _032_ _033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_37_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_87_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_204_ _014_ _017_ _018_ _019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_135_ _072_ _073_ _075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XANTENNA__250__A2 _033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_85_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
Xmacro_decap8_132 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_154 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_121 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_110 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_143 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmacro_decap8_187 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_176 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_165 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__150__A1 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XANTENNA__141__A1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_92_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XANTENNA__123__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_86_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_220_ _030_ _061_ net4 _032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_151_ net14 _091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_93_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_69_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_83_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_55_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_203_ net19 _018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_134_ _072_ _073_ _074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_93_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_0_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_80_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_66_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_47_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_62_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input20_I io_in[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmacro_decap8_111 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_100 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xmacro_decap8_133 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_155 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_144 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_122 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_53_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xmacro_decap8_188 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_177 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_166 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_90_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_44_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__227__I _116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_53_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_41_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_91_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_86_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_23_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_64_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_150_ net20 _087_ _090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_46_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
X_133_ _067_ net19 net6 _073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_202_ _015_ _016_ _017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_40_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_90_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_16
XFILLER_71_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_89_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xmacro_decap8_134 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_101 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_112 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_123 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
Xmacro_decap8_156 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA_input13_I io_in[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xmacro_decap8_145 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
Xmacro_decap8_189 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_178 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_167 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input5_I io_in[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_81_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_17_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_86_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_9_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_92_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_64_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
X_201_ _072_ _002_ _016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_132_ net7 _072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XANTENNA__161__I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XANTENNA__171__A1 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_32
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XFILLER_0_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XANTENNA__156__I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XANTENNA__153__A1 _090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
Xmacro_decap8_135 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_157 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_124 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_113 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_102 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xmacro_decap8_146 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
Xmacro_decap8_168 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
Xmacro_decap8_179 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_0_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XANTENNA__126__A1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_4
Xoutput30 net30 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_64
XFILLER_86_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
.ends

