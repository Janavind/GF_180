magic
tech gf180mcuC
magscale 1 10
timestamp 1670290001
<< metal1 >>
rect 74162 77198 74174 77250
rect 74226 77247 74238 77250
rect 75282 77247 75294 77250
rect 74226 77201 75294 77247
rect 74226 77198 74238 77201
rect 75282 77198 75294 77201
rect 75346 77198 75358 77250
rect 32386 76974 32398 77026
rect 32450 77023 32462 77026
rect 33282 77023 33294 77026
rect 32450 76977 33294 77023
rect 32450 76974 32462 76977
rect 33282 76974 33294 76977
rect 33346 76974 33358 77026
rect 37874 76974 37886 77026
rect 37938 77023 37950 77026
rect 38770 77023 38782 77026
rect 37938 76977 38782 77023
rect 37938 76974 37950 76977
rect 38770 76974 38782 76977
rect 38834 76974 38846 77026
rect 45378 76974 45390 77026
rect 45442 77023 45454 77026
rect 46722 77023 46734 77026
rect 45442 76977 46734 77023
rect 45442 76974 45454 76977
rect 46722 76974 46734 76977
rect 46786 76974 46798 77026
rect 48066 76974 48078 77026
rect 48130 77023 48142 77026
rect 48626 77023 48638 77026
rect 48130 76977 48638 77023
rect 48130 76974 48142 76977
rect 48626 76974 48638 76977
rect 48690 76974 48702 77026
rect 60722 76974 60734 77026
rect 60786 77023 60798 77026
rect 61282 77023 61294 77026
rect 60786 76977 61294 77023
rect 60786 76974 60798 76977
rect 61282 76974 61294 76977
rect 61346 76974 61358 77026
rect 76178 76974 76190 77026
rect 76242 77023 76254 77026
rect 76962 77023 76974 77026
rect 76242 76977 76974 77023
rect 76242 76974 76254 76977
rect 76962 76974 76974 76977
rect 77026 76974 77038 77026
rect 1344 76858 78624 76892
rect 1344 76806 19838 76858
rect 19890 76806 19942 76858
rect 19994 76806 20046 76858
rect 20098 76806 50558 76858
rect 50610 76806 50662 76858
rect 50714 76806 50766 76858
rect 50818 76806 78624 76858
rect 1344 76772 78624 76806
rect 3838 76690 3890 76702
rect 3838 76626 3890 76638
rect 4958 76690 5010 76702
rect 4958 76626 5010 76638
rect 7870 76690 7922 76702
rect 7870 76626 7922 76638
rect 8878 76690 8930 76702
rect 8878 76626 8930 76638
rect 9886 76690 9938 76702
rect 9886 76626 9938 76638
rect 11006 76690 11058 76702
rect 11006 76626 11058 76638
rect 43374 76690 43426 76702
rect 47070 76690 47122 76702
rect 55806 76690 55858 76702
rect 46722 76638 46734 76690
rect 46786 76638 46798 76690
rect 51650 76638 51662 76690
rect 51714 76638 51726 76690
rect 43374 76626 43426 76638
rect 47070 76626 47122 76638
rect 55806 76626 55858 76638
rect 61294 76690 61346 76702
rect 61294 76626 61346 76638
rect 61854 76690 61906 76702
rect 61854 76626 61906 76638
rect 62526 76690 62578 76702
rect 62526 76626 62578 76638
rect 63198 76690 63250 76702
rect 63198 76626 63250 76638
rect 72382 76690 72434 76702
rect 72382 76626 72434 76638
rect 73054 76690 73106 76702
rect 73054 76626 73106 76638
rect 73950 76690 74002 76702
rect 73950 76626 74002 76638
rect 74622 76690 74674 76702
rect 74622 76626 74674 76638
rect 75294 76690 75346 76702
rect 75294 76626 75346 76638
rect 76302 76690 76354 76702
rect 76302 76626 76354 76638
rect 76974 76690 77026 76702
rect 76974 76626 77026 76638
rect 77758 76690 77810 76702
rect 77758 76626 77810 76638
rect 29486 76578 29538 76590
rect 32398 76578 32450 76590
rect 1922 76526 1934 76578
rect 1986 76526 1998 76578
rect 5842 76526 5854 76578
rect 5906 76526 5918 76578
rect 11666 76526 11678 76578
rect 11730 76526 11742 76578
rect 13794 76526 13806 76578
rect 13858 76526 13870 76578
rect 17714 76526 17726 76578
rect 17778 76526 17790 76578
rect 30146 76526 30158 76578
rect 30210 76526 30222 76578
rect 29486 76514 29538 76526
rect 32398 76514 32450 76526
rect 37214 76578 37266 76590
rect 37214 76514 37266 76526
rect 38110 76578 38162 76590
rect 44942 76578 44994 76590
rect 38882 76526 38894 76578
rect 38946 76526 38958 76578
rect 42018 76526 42030 76578
rect 42082 76526 42094 76578
rect 38110 76514 38162 76526
rect 44942 76514 44994 76526
rect 45278 76578 45330 76590
rect 45278 76514 45330 76526
rect 45838 76578 45890 76590
rect 45838 76514 45890 76526
rect 47742 76578 47794 76590
rect 47742 76514 47794 76526
rect 48078 76578 48130 76590
rect 48078 76514 48130 76526
rect 48974 76578 49026 76590
rect 48974 76514 49026 76526
rect 49870 76578 49922 76590
rect 49870 76514 49922 76526
rect 50094 76578 50146 76590
rect 50094 76514 50146 76526
rect 50766 76578 50818 76590
rect 50766 76514 50818 76526
rect 50990 76578 51042 76590
rect 58942 76578 58994 76590
rect 54786 76526 54798 76578
rect 54850 76526 54862 76578
rect 57922 76526 57934 76578
rect 57986 76526 57998 76578
rect 50990 76514 51042 76526
rect 58942 76514 58994 76526
rect 59278 76578 59330 76590
rect 64430 76578 64482 76590
rect 71486 76578 71538 76590
rect 60946 76526 60958 76578
rect 61010 76526 61022 76578
rect 67218 76526 67230 76578
rect 67282 76526 67294 76578
rect 70578 76526 70590 76578
rect 70642 76526 70654 76578
rect 59278 76514 59330 76526
rect 64430 76514 64482 76526
rect 71486 76514 71538 76526
rect 37102 76466 37154 76478
rect 43262 76466 43314 76478
rect 6850 76414 6862 76466
rect 6914 76414 6926 76466
rect 12786 76414 12798 76466
rect 12850 76414 12862 76466
rect 14914 76414 14926 76466
rect 14978 76414 14990 76466
rect 16706 76414 16718 76466
rect 16770 76414 16782 76466
rect 18834 76414 18846 76466
rect 18898 76414 18910 76466
rect 20626 76414 20638 76466
rect 20690 76414 20702 76466
rect 22754 76414 22766 76466
rect 22818 76414 22830 76466
rect 24546 76414 24558 76466
rect 24610 76414 24622 76466
rect 26562 76414 26574 76466
rect 26626 76414 26638 76466
rect 28466 76414 28478 76466
rect 28530 76414 28542 76466
rect 31042 76414 31054 76466
rect 31106 76414 31118 76466
rect 32162 76414 32174 76466
rect 32226 76414 32238 76466
rect 33282 76414 33294 76466
rect 33346 76414 33358 76466
rect 35074 76414 35086 76466
rect 35138 76414 35150 76466
rect 43026 76414 43038 76466
rect 43090 76414 43102 76466
rect 37102 76402 37154 76414
rect 43262 76402 43314 76414
rect 43486 76466 43538 76478
rect 43486 76402 43538 76414
rect 43598 76466 43650 76478
rect 43598 76402 43650 76414
rect 46174 76466 46226 76478
rect 46174 76402 46226 76414
rect 49086 76466 49138 76478
rect 51102 76466 51154 76478
rect 49634 76414 49646 76466
rect 49698 76414 49710 76466
rect 49086 76402 49138 76414
rect 51102 76402 51154 76414
rect 51998 76466 52050 76478
rect 51998 76402 52050 76414
rect 63758 76466 63810 76478
rect 73266 76414 73278 76466
rect 73330 76414 73342 76466
rect 63758 76402 63810 76414
rect 37886 76354 37938 76366
rect 44270 76354 44322 76366
rect 59726 76354 59778 76366
rect 3266 76302 3278 76354
rect 3330 76302 3342 76354
rect 15698 76302 15710 76354
rect 15762 76302 15774 76354
rect 19618 76302 19630 76354
rect 19682 76302 19694 76354
rect 21858 76302 21870 76354
rect 21922 76302 21934 76354
rect 23762 76302 23774 76354
rect 23826 76302 23838 76354
rect 25778 76302 25790 76354
rect 25842 76302 25854 76354
rect 27794 76302 27806 76354
rect 27858 76302 27870 76354
rect 33954 76302 33966 76354
rect 34018 76302 34030 76354
rect 35858 76302 35870 76354
rect 35922 76302 35934 76354
rect 40226 76302 40238 76354
rect 40290 76302 40302 76354
rect 41010 76302 41022 76354
rect 41074 76302 41086 76354
rect 49970 76302 49982 76354
rect 50034 76302 50046 76354
rect 56914 76302 56926 76354
rect 56978 76302 56990 76354
rect 37886 76290 37938 76302
rect 44270 76290 44322 76302
rect 59726 76290 59778 76302
rect 37214 76242 37266 76254
rect 37214 76178 37266 76190
rect 38222 76242 38274 76254
rect 38222 76178 38274 76190
rect 48974 76242 49026 76254
rect 48974 76178 49026 76190
rect 52670 76242 52722 76254
rect 52670 76178 52722 76190
rect 64878 76242 64930 76254
rect 64878 76178 64930 76190
rect 68350 76242 68402 76254
rect 68350 76178 68402 76190
rect 1344 76074 78624 76108
rect 1344 76022 4478 76074
rect 4530 76022 4582 76074
rect 4634 76022 4686 76074
rect 4738 76022 35198 76074
rect 35250 76022 35302 76074
rect 35354 76022 35406 76074
rect 35458 76022 65918 76074
rect 65970 76022 66022 76074
rect 66074 76022 66126 76074
rect 66178 76022 78624 76074
rect 1344 75988 78624 76022
rect 46734 75906 46786 75918
rect 37874 75903 37886 75906
rect 37329 75857 37886 75903
rect 1822 75794 1874 75806
rect 1822 75730 1874 75742
rect 7870 75794 7922 75806
rect 7870 75730 7922 75742
rect 19854 75794 19906 75806
rect 19854 75730 19906 75742
rect 20862 75794 20914 75806
rect 20862 75730 20914 75742
rect 23998 75794 24050 75806
rect 23998 75730 24050 75742
rect 24782 75794 24834 75806
rect 32722 75742 32734 75794
rect 32786 75742 32798 75794
rect 36194 75742 36206 75794
rect 36258 75742 36270 75794
rect 24782 75730 24834 75742
rect 12910 75682 12962 75694
rect 12910 75618 12962 75630
rect 15822 75682 15874 75694
rect 15822 75618 15874 75630
rect 17838 75682 17890 75694
rect 17838 75618 17890 75630
rect 26574 75682 26626 75694
rect 26574 75618 26626 75630
rect 30158 75682 30210 75694
rect 30158 75618 30210 75630
rect 30382 75682 30434 75694
rect 31278 75682 31330 75694
rect 30930 75630 30942 75682
rect 30994 75630 31006 75682
rect 30382 75618 30434 75630
rect 31278 75618 31330 75630
rect 31502 75682 31554 75694
rect 32050 75630 32062 75682
rect 32114 75630 32126 75682
rect 36082 75630 36094 75682
rect 36146 75630 36158 75682
rect 31502 75618 31554 75630
rect 5854 75570 5906 75582
rect 5854 75506 5906 75518
rect 7198 75570 7250 75582
rect 7198 75506 7250 75518
rect 13694 75570 13746 75582
rect 13694 75506 13746 75518
rect 15262 75570 15314 75582
rect 15262 75506 15314 75518
rect 17278 75570 17330 75582
rect 17278 75506 17330 75518
rect 19294 75570 19346 75582
rect 19294 75506 19346 75518
rect 21646 75570 21698 75582
rect 21646 75506 21698 75518
rect 23326 75570 23378 75582
rect 23326 75506 23378 75518
rect 25342 75570 25394 75582
rect 25342 75506 25394 75518
rect 27134 75570 27186 75582
rect 27134 75506 27186 75518
rect 27918 75570 27970 75582
rect 27918 75506 27970 75518
rect 28478 75570 28530 75582
rect 28478 75506 28530 75518
rect 28814 75570 28866 75582
rect 33854 75570 33906 75582
rect 29810 75518 29822 75570
rect 29874 75518 29886 75570
rect 28814 75506 28866 75518
rect 33854 75506 33906 75518
rect 34078 75570 34130 75582
rect 34078 75506 34130 75518
rect 34302 75570 34354 75582
rect 34302 75506 34354 75518
rect 34414 75570 34466 75582
rect 34414 75506 34466 75518
rect 35198 75570 35250 75582
rect 35198 75506 35250 75518
rect 35534 75570 35586 75582
rect 35534 75506 35586 75518
rect 36766 75570 36818 75582
rect 36766 75506 36818 75518
rect 36318 75458 36370 75470
rect 36318 75394 36370 75406
rect 36542 75458 36594 75470
rect 37329 75458 37375 75857
rect 37874 75854 37886 75857
rect 37938 75854 37950 75906
rect 40898 75854 40910 75906
rect 40962 75903 40974 75906
rect 41570 75903 41582 75906
rect 40962 75857 41582 75903
rect 40962 75854 40974 75857
rect 41570 75854 41582 75857
rect 41634 75854 41646 75906
rect 43474 75854 43486 75906
rect 43538 75854 43550 75906
rect 46734 75842 46786 75854
rect 57262 75906 57314 75918
rect 57262 75842 57314 75854
rect 70926 75906 70978 75918
rect 70926 75842 70978 75854
rect 40462 75794 40514 75806
rect 38770 75742 38782 75794
rect 38834 75742 38846 75794
rect 40462 75730 40514 75742
rect 46286 75794 46338 75806
rect 46286 75730 46338 75742
rect 49758 75794 49810 75806
rect 49758 75730 49810 75742
rect 50878 75794 50930 75806
rect 50878 75730 50930 75742
rect 52558 75794 52610 75806
rect 52558 75730 52610 75742
rect 54126 75794 54178 75806
rect 62862 75794 62914 75806
rect 56354 75742 56366 75794
rect 56418 75742 56430 75794
rect 56914 75742 56926 75794
rect 56978 75742 56990 75794
rect 54126 75730 54178 75742
rect 62862 75730 62914 75742
rect 68686 75794 68738 75806
rect 68686 75730 68738 75742
rect 40686 75682 40738 75694
rect 38098 75630 38110 75682
rect 38162 75630 38174 75682
rect 40686 75618 40738 75630
rect 43038 75682 43090 75694
rect 43038 75618 43090 75630
rect 50766 75682 50818 75694
rect 50766 75618 50818 75630
rect 50990 75682 51042 75694
rect 50990 75618 51042 75630
rect 51774 75682 51826 75694
rect 51774 75618 51826 75630
rect 52222 75682 52274 75694
rect 52222 75618 52274 75630
rect 54350 75682 54402 75694
rect 54350 75618 54402 75630
rect 61294 75682 61346 75694
rect 61294 75618 61346 75630
rect 61630 75682 61682 75694
rect 61630 75618 61682 75630
rect 62190 75682 62242 75694
rect 62190 75618 62242 75630
rect 73950 75682 74002 75694
rect 73950 75618 74002 75630
rect 40014 75570 40066 75582
rect 40014 75506 40066 75518
rect 41806 75570 41858 75582
rect 41806 75506 41858 75518
rect 42814 75570 42866 75582
rect 42814 75506 42866 75518
rect 42926 75570 42978 75582
rect 42926 75506 42978 75518
rect 44382 75570 44434 75582
rect 44382 75506 44434 75518
rect 45838 75570 45890 75582
rect 53678 75570 53730 75582
rect 58158 75570 58210 75582
rect 48850 75518 48862 75570
rect 48914 75518 48926 75570
rect 55010 75518 55022 75570
rect 55074 75518 55086 75570
rect 45838 75506 45890 75518
rect 53678 75506 53730 75518
rect 58158 75506 58210 75518
rect 59950 75570 60002 75582
rect 59950 75506 60002 75518
rect 60510 75570 60562 75582
rect 60510 75506 60562 75518
rect 62302 75570 62354 75582
rect 66670 75570 66722 75582
rect 64978 75518 64990 75570
rect 65042 75518 65054 75570
rect 62302 75506 62354 75518
rect 66670 75506 66722 75518
rect 68014 75570 68066 75582
rect 70254 75570 70306 75582
rect 77198 75570 77250 75582
rect 69346 75518 69358 75570
rect 69410 75518 69422 75570
rect 73042 75518 73054 75570
rect 73106 75518 73118 75570
rect 76066 75518 76078 75570
rect 76130 75518 76142 75570
rect 68014 75506 68066 75518
rect 70254 75506 70306 75518
rect 77198 75506 77250 75518
rect 78094 75570 78146 75582
rect 78094 75506 78146 75518
rect 37662 75458 37714 75470
rect 37314 75406 37326 75458
rect 37378 75406 37390 75458
rect 36542 75394 36594 75406
rect 37662 75394 37714 75406
rect 40126 75458 40178 75470
rect 40126 75394 40178 75406
rect 40238 75458 40290 75470
rect 40238 75394 40290 75406
rect 41246 75458 41298 75470
rect 41246 75394 41298 75406
rect 42142 75458 42194 75470
rect 42142 75394 42194 75406
rect 44046 75458 44098 75470
rect 44046 75394 44098 75406
rect 45502 75458 45554 75470
rect 45502 75394 45554 75406
rect 50542 75458 50594 75470
rect 50542 75394 50594 75406
rect 51550 75458 51602 75470
rect 51550 75394 51602 75406
rect 51662 75458 51714 75470
rect 51662 75394 51714 75406
rect 53790 75458 53842 75470
rect 53790 75394 53842 75406
rect 53902 75458 53954 75470
rect 53902 75394 53954 75406
rect 57038 75458 57090 75470
rect 57038 75394 57090 75406
rect 57822 75458 57874 75470
rect 59054 75458 59106 75470
rect 58706 75406 58718 75458
rect 58770 75406 58782 75458
rect 57822 75394 57874 75406
rect 59054 75394 59106 75406
rect 59614 75458 59666 75470
rect 59614 75394 59666 75406
rect 61518 75458 61570 75470
rect 61518 75394 61570 75406
rect 65998 75458 66050 75470
rect 65998 75394 66050 75406
rect 67342 75458 67394 75470
rect 67342 75394 67394 75406
rect 69694 75458 69746 75470
rect 69694 75394 69746 75406
rect 1344 75290 78624 75324
rect 1344 75238 19838 75290
rect 19890 75238 19942 75290
rect 19994 75238 20046 75290
rect 20098 75238 50558 75290
rect 50610 75238 50662 75290
rect 50714 75238 50766 75290
rect 50818 75238 78624 75290
rect 1344 75204 78624 75238
rect 28142 75122 28194 75134
rect 28142 75058 28194 75070
rect 29038 75122 29090 75134
rect 29038 75058 29090 75070
rect 30270 75122 30322 75134
rect 30270 75058 30322 75070
rect 30942 75122 30994 75134
rect 34302 75122 34354 75134
rect 36542 75122 36594 75134
rect 32274 75070 32286 75122
rect 32338 75070 32350 75122
rect 35298 75070 35310 75122
rect 35362 75070 35374 75122
rect 30942 75058 30994 75070
rect 34302 75058 34354 75070
rect 36542 75058 36594 75070
rect 39454 75122 39506 75134
rect 39454 75058 39506 75070
rect 39678 75122 39730 75134
rect 39678 75058 39730 75070
rect 39790 75122 39842 75134
rect 39790 75058 39842 75070
rect 40798 75122 40850 75134
rect 40798 75058 40850 75070
rect 41694 75122 41746 75134
rect 41694 75058 41746 75070
rect 41806 75122 41858 75134
rect 41806 75058 41858 75070
rect 44270 75122 44322 75134
rect 46734 75122 46786 75134
rect 44706 75070 44718 75122
rect 44770 75070 44782 75122
rect 44270 75058 44322 75070
rect 46734 75058 46786 75070
rect 47518 75122 47570 75134
rect 47518 75058 47570 75070
rect 50094 75122 50146 75134
rect 55358 75122 55410 75134
rect 54226 75070 54238 75122
rect 54290 75070 54302 75122
rect 50094 75058 50146 75070
rect 55358 75058 55410 75070
rect 57598 75122 57650 75134
rect 57598 75058 57650 75070
rect 60622 75122 60674 75134
rect 60622 75058 60674 75070
rect 61966 75122 62018 75134
rect 61966 75058 62018 75070
rect 62638 75122 62690 75134
rect 62638 75058 62690 75070
rect 63310 75122 63362 75134
rect 63310 75058 63362 75070
rect 63982 75122 64034 75134
rect 63982 75058 64034 75070
rect 65438 75122 65490 75134
rect 65438 75058 65490 75070
rect 68350 75122 68402 75134
rect 68350 75058 68402 75070
rect 69134 75122 69186 75134
rect 69134 75058 69186 75070
rect 70814 75122 70866 75134
rect 70814 75058 70866 75070
rect 73278 75122 73330 75134
rect 73278 75058 73330 75070
rect 31166 75010 31218 75022
rect 31166 74946 31218 74958
rect 33742 75010 33794 75022
rect 38782 75010 38834 75022
rect 45502 75010 45554 75022
rect 37426 74958 37438 75010
rect 37490 74958 37502 75010
rect 40450 74958 40462 75010
rect 40514 74958 40526 75010
rect 33742 74946 33794 74958
rect 38782 74946 38834 74958
rect 45502 74946 45554 74958
rect 46846 75010 46898 75022
rect 49982 75010 50034 75022
rect 48626 74958 48638 75010
rect 48690 74958 48702 75010
rect 46846 74946 46898 74958
rect 49982 74946 50034 74958
rect 50318 75010 50370 75022
rect 50318 74946 50370 74958
rect 53006 75010 53058 75022
rect 55246 75010 55298 75022
rect 54114 74958 54126 75010
rect 54178 74958 54190 75010
rect 53006 74946 53058 74958
rect 55246 74946 55298 74958
rect 56366 75010 56418 75022
rect 56366 74946 56418 74958
rect 56702 75010 56754 75022
rect 60734 75010 60786 75022
rect 58146 74958 58158 75010
rect 58210 74958 58222 75010
rect 58706 74958 58718 75010
rect 58770 74958 58782 75010
rect 77634 74958 77646 75010
rect 77698 74958 77710 75010
rect 56702 74946 56754 74958
rect 60734 74946 60786 74958
rect 29374 74898 29426 74910
rect 30718 74898 30770 74910
rect 30034 74846 30046 74898
rect 30098 74846 30110 74898
rect 29374 74834 29426 74846
rect 30718 74834 30770 74846
rect 31278 74898 31330 74910
rect 31278 74834 31330 74846
rect 32846 74898 32898 74910
rect 32846 74834 32898 74846
rect 34190 74898 34242 74910
rect 34190 74834 34242 74846
rect 34526 74898 34578 74910
rect 34526 74834 34578 74846
rect 34638 74898 34690 74910
rect 38446 74898 38498 74910
rect 37650 74846 37662 74898
rect 37714 74846 37726 74898
rect 34638 74834 34690 74846
rect 38446 74834 38498 74846
rect 39902 74898 39954 74910
rect 39902 74834 39954 74846
rect 41582 74898 41634 74910
rect 41582 74834 41634 74846
rect 42702 74898 42754 74910
rect 44158 74898 44210 74910
rect 42914 74846 42926 74898
rect 42978 74846 42990 74898
rect 43474 74846 43486 74898
rect 43538 74846 43550 74898
rect 42702 74834 42754 74846
rect 44158 74834 44210 74846
rect 44494 74898 44546 74910
rect 44494 74834 44546 74846
rect 44718 74898 44770 74910
rect 44718 74834 44770 74846
rect 45726 74898 45778 74910
rect 45726 74834 45778 74846
rect 46174 74898 46226 74910
rect 46174 74834 46226 74846
rect 46510 74898 46562 74910
rect 46510 74834 46562 74846
rect 47854 74898 47906 74910
rect 53902 74898 53954 74910
rect 48514 74846 48526 74898
rect 48578 74846 48590 74898
rect 49522 74846 49534 74898
rect 49586 74846 49598 74898
rect 51650 74846 51662 74898
rect 51714 74846 51726 74898
rect 53218 74846 53230 74898
rect 53282 74846 53294 74898
rect 47854 74834 47906 74846
rect 53902 74834 53954 74846
rect 54350 74898 54402 74910
rect 55470 74898 55522 74910
rect 54674 74846 54686 74898
rect 54738 74846 54750 74898
rect 54350 74834 54402 74846
rect 55470 74834 55522 74846
rect 55918 74898 55970 74910
rect 55918 74834 55970 74846
rect 59390 74898 59442 74910
rect 59390 74834 59442 74846
rect 59614 74898 59666 74910
rect 61406 74898 61458 74910
rect 59938 74846 59950 74898
rect 60002 74846 60014 74898
rect 59614 74834 59666 74846
rect 61406 74834 61458 74846
rect 28590 74786 28642 74798
rect 28590 74722 28642 74734
rect 32622 74786 32674 74798
rect 32622 74722 32674 74734
rect 35870 74786 35922 74798
rect 35870 74722 35922 74734
rect 42814 74786 42866 74798
rect 42814 74722 42866 74734
rect 45614 74786 45666 74798
rect 51214 74786 51266 74798
rect 59502 74786 59554 74798
rect 49970 74734 49982 74786
rect 50034 74734 50046 74786
rect 52098 74734 52110 74786
rect 52162 74734 52174 74786
rect 45614 74722 45666 74734
rect 51214 74722 51266 74734
rect 59502 74722 59554 74734
rect 64542 74786 64594 74798
rect 64542 74722 64594 74734
rect 35646 74674 35698 74686
rect 35646 74610 35698 74622
rect 36878 74674 36930 74686
rect 57934 74674 57986 74686
rect 43250 74622 43262 74674
rect 43314 74622 43326 74674
rect 36878 74610 36930 74622
rect 57934 74610 57986 74622
rect 60622 74674 60674 74686
rect 60622 74610 60674 74622
rect 61294 74674 61346 74686
rect 61294 74610 61346 74622
rect 74510 74674 74562 74686
rect 74510 74610 74562 74622
rect 1344 74506 78624 74540
rect 1344 74454 4478 74506
rect 4530 74454 4582 74506
rect 4634 74454 4686 74506
rect 4738 74454 35198 74506
rect 35250 74454 35302 74506
rect 35354 74454 35406 74506
rect 35458 74454 65918 74506
rect 65970 74454 66022 74506
rect 66074 74454 66126 74506
rect 66178 74454 78624 74506
rect 1344 74420 78624 74454
rect 32286 74338 32338 74350
rect 32286 74274 32338 74286
rect 33070 74338 33122 74350
rect 44270 74338 44322 74350
rect 34178 74286 34190 74338
rect 34242 74286 34254 74338
rect 33070 74274 33122 74286
rect 44270 74274 44322 74286
rect 44382 74338 44434 74350
rect 44382 74274 44434 74286
rect 45726 74338 45778 74350
rect 45726 74274 45778 74286
rect 48414 74338 48466 74350
rect 51662 74338 51714 74350
rect 49746 74286 49758 74338
rect 49810 74286 49822 74338
rect 48414 74274 48466 74286
rect 51662 74274 51714 74286
rect 56142 74338 56194 74350
rect 56142 74274 56194 74286
rect 57038 74338 57090 74350
rect 57038 74274 57090 74286
rect 59838 74338 59890 74350
rect 59838 74274 59890 74286
rect 28814 74226 28866 74238
rect 28814 74162 28866 74174
rect 29710 74226 29762 74238
rect 29710 74162 29762 74174
rect 32174 74226 32226 74238
rect 32174 74162 32226 74174
rect 32846 74226 32898 74238
rect 32846 74162 32898 74174
rect 34526 74226 34578 74238
rect 40126 74226 40178 74238
rect 44046 74226 44098 74238
rect 37986 74174 37998 74226
rect 38050 74174 38062 74226
rect 42130 74174 42142 74226
rect 42194 74174 42206 74226
rect 42690 74174 42702 74226
rect 42754 74174 42766 74226
rect 34526 74162 34578 74174
rect 40126 74162 40178 74174
rect 44046 74162 44098 74174
rect 45950 74226 46002 74238
rect 45950 74162 46002 74174
rect 48526 74226 48578 74238
rect 54238 74226 54290 74238
rect 54002 74174 54014 74226
rect 54066 74174 54078 74226
rect 48526 74162 48578 74174
rect 54238 74162 54290 74174
rect 56366 74226 56418 74238
rect 61966 74226 62018 74238
rect 57362 74174 57374 74226
rect 57426 74174 57438 74226
rect 56366 74162 56418 74174
rect 61966 74162 62018 74174
rect 62414 74226 62466 74238
rect 62414 74162 62466 74174
rect 62862 74226 62914 74238
rect 62862 74162 62914 74174
rect 63310 74226 63362 74238
rect 63310 74162 63362 74174
rect 78094 74226 78146 74238
rect 78094 74162 78146 74174
rect 34750 74114 34802 74126
rect 31938 74062 31950 74114
rect 32002 74062 32014 74114
rect 34750 74050 34802 74062
rect 35310 74114 35362 74126
rect 35310 74050 35362 74062
rect 35534 74114 35586 74126
rect 35534 74050 35586 74062
rect 35982 74114 36034 74126
rect 35982 74050 36034 74062
rect 36542 74114 36594 74126
rect 36542 74050 36594 74062
rect 36878 74114 36930 74126
rect 38894 74114 38946 74126
rect 37538 74062 37550 74114
rect 37602 74062 37614 74114
rect 36878 74050 36930 74062
rect 38894 74050 38946 74062
rect 39566 74114 39618 74126
rect 39566 74050 39618 74062
rect 40574 74114 40626 74126
rect 40574 74050 40626 74062
rect 40686 74114 40738 74126
rect 40686 74050 40738 74062
rect 40798 74114 40850 74126
rect 40798 74050 40850 74062
rect 41246 74114 41298 74126
rect 43934 74114 43986 74126
rect 42018 74062 42030 74114
rect 42082 74062 42094 74114
rect 43026 74062 43038 74114
rect 43090 74062 43102 74114
rect 41246 74050 41298 74062
rect 43934 74050 43986 74062
rect 46174 74114 46226 74126
rect 46174 74050 46226 74062
rect 46398 74114 46450 74126
rect 51102 74114 51154 74126
rect 50530 74062 50542 74114
rect 50594 74062 50606 74114
rect 46398 74050 46450 74062
rect 51102 74050 51154 74062
rect 52222 74114 52274 74126
rect 52222 74050 52274 74062
rect 52558 74114 52610 74126
rect 55470 74114 55522 74126
rect 53442 74062 53454 74114
rect 53506 74062 53518 74114
rect 54450 74062 54462 74114
rect 54514 74062 54526 74114
rect 52558 74050 52610 74062
rect 55470 74050 55522 74062
rect 55918 74114 55970 74126
rect 55918 74050 55970 74062
rect 59166 74114 59218 74126
rect 59166 74050 59218 74062
rect 59390 74114 59442 74126
rect 59390 74050 59442 74062
rect 59614 74114 59666 74126
rect 59614 74050 59666 74062
rect 60286 74114 60338 74126
rect 60286 74050 60338 74062
rect 30158 74002 30210 74014
rect 30158 73938 30210 73950
rect 30494 74002 30546 74014
rect 30494 73938 30546 73950
rect 31054 74002 31106 74014
rect 31054 73938 31106 73950
rect 35422 74002 35474 74014
rect 35422 73938 35474 73950
rect 37998 74002 38050 74014
rect 37998 73938 38050 73950
rect 38110 74002 38162 74014
rect 38110 73938 38162 73950
rect 39006 74002 39058 74014
rect 50206 74002 50258 74014
rect 42242 73950 42254 74002
rect 42306 73950 42318 74002
rect 39006 73938 39058 73950
rect 50206 73938 50258 73950
rect 50318 74002 50370 74014
rect 50318 73938 50370 73950
rect 51326 74002 51378 74014
rect 51326 73938 51378 73950
rect 51774 74002 51826 74014
rect 57262 74002 57314 74014
rect 53554 73950 53566 74002
rect 53618 73950 53630 74002
rect 51774 73938 51826 73950
rect 57262 73938 57314 73950
rect 57934 74002 57986 74014
rect 57934 73938 57986 73950
rect 58270 74002 58322 74014
rect 58270 73938 58322 73950
rect 60622 74002 60674 74014
rect 60622 73938 60674 73950
rect 31390 73890 31442 73902
rect 36654 73890 36706 73902
rect 33394 73838 33406 73890
rect 33458 73838 33470 73890
rect 31390 73826 31442 73838
rect 36654 73826 36706 73838
rect 38334 73890 38386 73902
rect 38334 73826 38386 73838
rect 39118 73890 39170 73902
rect 39118 73826 39170 73838
rect 46286 73890 46338 73902
rect 46286 73826 46338 73838
rect 47070 73890 47122 73902
rect 47070 73826 47122 73838
rect 47742 73890 47794 73902
rect 47742 73826 47794 73838
rect 49086 73890 49138 73902
rect 49086 73826 49138 73838
rect 51550 73890 51602 73902
rect 51550 73826 51602 73838
rect 52446 73890 52498 73902
rect 52446 73826 52498 73838
rect 58046 73890 58098 73902
rect 58046 73826 58098 73838
rect 59278 73890 59330 73902
rect 59278 73826 59330 73838
rect 60510 73890 60562 73902
rect 60510 73826 60562 73838
rect 61406 73890 61458 73902
rect 61406 73826 61458 73838
rect 1344 73722 78624 73756
rect 1344 73670 19838 73722
rect 19890 73670 19942 73722
rect 19994 73670 20046 73722
rect 20098 73670 50558 73722
rect 50610 73670 50662 73722
rect 50714 73670 50766 73722
rect 50818 73670 78624 73722
rect 1344 73636 78624 73670
rect 29486 73554 29538 73566
rect 29486 73490 29538 73502
rect 30494 73554 30546 73566
rect 30494 73490 30546 73502
rect 31390 73554 31442 73566
rect 31390 73490 31442 73502
rect 32062 73554 32114 73566
rect 32062 73490 32114 73502
rect 32958 73554 33010 73566
rect 32958 73490 33010 73502
rect 33630 73554 33682 73566
rect 33630 73490 33682 73502
rect 34862 73554 34914 73566
rect 34862 73490 34914 73502
rect 35758 73554 35810 73566
rect 35758 73490 35810 73502
rect 36430 73554 36482 73566
rect 36430 73490 36482 73502
rect 40238 73554 40290 73566
rect 40238 73490 40290 73502
rect 40350 73554 40402 73566
rect 40350 73490 40402 73502
rect 40574 73554 40626 73566
rect 40574 73490 40626 73502
rect 41470 73554 41522 73566
rect 41470 73490 41522 73502
rect 41694 73554 41746 73566
rect 41694 73490 41746 73502
rect 43822 73554 43874 73566
rect 43822 73490 43874 73502
rect 47518 73554 47570 73566
rect 47518 73490 47570 73502
rect 50542 73554 50594 73566
rect 50542 73490 50594 73502
rect 55470 73554 55522 73566
rect 55470 73490 55522 73502
rect 56142 73554 56194 73566
rect 56142 73490 56194 73502
rect 56254 73554 56306 73566
rect 56254 73490 56306 73502
rect 57598 73554 57650 73566
rect 57598 73490 57650 73502
rect 60846 73554 60898 73566
rect 60846 73490 60898 73502
rect 61406 73554 61458 73566
rect 61406 73490 61458 73502
rect 61854 73554 61906 73566
rect 61854 73490 61906 73502
rect 62302 73554 62354 73566
rect 62302 73490 62354 73502
rect 62862 73554 62914 73566
rect 62862 73490 62914 73502
rect 31278 73442 31330 73454
rect 31278 73378 31330 73390
rect 31502 73442 31554 73454
rect 31502 73378 31554 73390
rect 34526 73442 34578 73454
rect 40798 73442 40850 73454
rect 37538 73390 37550 73442
rect 37602 73390 37614 73442
rect 34526 73378 34578 73390
rect 40798 73378 40850 73390
rect 41806 73442 41858 73454
rect 41806 73378 41858 73390
rect 45390 73442 45442 73454
rect 45390 73378 45442 73390
rect 48526 73442 48578 73454
rect 48526 73378 48578 73390
rect 48750 73442 48802 73454
rect 48750 73378 48802 73390
rect 51102 73442 51154 73454
rect 54462 73442 54514 73454
rect 51762 73390 51774 73442
rect 51826 73390 51838 73442
rect 52770 73390 52782 73442
rect 52834 73390 52846 73442
rect 51102 73378 51154 73390
rect 54462 73378 54514 73390
rect 57822 73442 57874 73454
rect 57822 73378 57874 73390
rect 60286 73442 60338 73454
rect 60286 73378 60338 73390
rect 38222 73330 38274 73342
rect 44606 73330 44658 73342
rect 33842 73278 33854 73330
rect 33906 73278 33918 73330
rect 37426 73278 37438 73330
rect 37490 73278 37502 73330
rect 38658 73278 38670 73330
rect 38722 73278 38734 73330
rect 38222 73266 38274 73278
rect 44606 73266 44658 73278
rect 45278 73330 45330 73342
rect 54574 73330 54626 73342
rect 46386 73278 46398 73330
rect 46450 73278 46462 73330
rect 51874 73278 51886 73330
rect 51938 73278 51950 73330
rect 52546 73278 52558 73330
rect 52610 73278 52622 73330
rect 53554 73278 53566 73330
rect 53618 73278 53630 73330
rect 45278 73266 45330 73278
rect 54574 73266 54626 73278
rect 54798 73330 54850 73342
rect 54798 73266 54850 73278
rect 56030 73330 56082 73342
rect 56030 73266 56082 73278
rect 56702 73330 56754 73342
rect 59042 73278 59054 73330
rect 59106 73278 59118 73330
rect 56702 73266 56754 73278
rect 29934 73218 29986 73230
rect 29934 73154 29986 73166
rect 30382 73218 30434 73230
rect 39790 73218 39842 73230
rect 39106 73166 39118 73218
rect 39170 73166 39182 73218
rect 30382 73154 30434 73166
rect 39790 73154 39842 73166
rect 42590 73218 42642 73230
rect 42590 73154 42642 73166
rect 45950 73218 46002 73230
rect 48638 73218 48690 73230
rect 46274 73166 46286 73218
rect 46338 73166 46350 73218
rect 45950 73154 46002 73166
rect 48638 73154 48690 73166
rect 49646 73218 49698 73230
rect 58606 73218 58658 73230
rect 52098 73166 52110 73218
rect 52162 73166 52174 73218
rect 59378 73166 59390 73218
rect 59442 73166 59454 73218
rect 49646 73154 49698 73166
rect 58606 73154 58658 73166
rect 36766 73106 36818 73118
rect 36766 73042 36818 73054
rect 42814 73106 42866 73118
rect 42814 73042 42866 73054
rect 43038 73106 43090 73118
rect 43038 73042 43090 73054
rect 43486 73106 43538 73118
rect 43486 73042 43538 73054
rect 44830 73106 44882 73118
rect 44830 73042 44882 73054
rect 45278 73106 45330 73118
rect 45278 73042 45330 73054
rect 49870 73106 49922 73118
rect 49870 73042 49922 73054
rect 50094 73106 50146 73118
rect 50094 73042 50146 73054
rect 50990 73106 51042 73118
rect 50990 73042 51042 73054
rect 54910 73106 54962 73118
rect 54910 73042 54962 73054
rect 57486 73106 57538 73118
rect 57486 73042 57538 73054
rect 60174 73106 60226 73118
rect 60174 73042 60226 73054
rect 1344 72938 78624 72972
rect 1344 72886 4478 72938
rect 4530 72886 4582 72938
rect 4634 72886 4686 72938
rect 4738 72886 35198 72938
rect 35250 72886 35302 72938
rect 35354 72886 35406 72938
rect 35458 72886 65918 72938
rect 65970 72886 66022 72938
rect 66074 72886 66126 72938
rect 66178 72886 78624 72938
rect 1344 72852 78624 72886
rect 36654 72770 36706 72782
rect 36654 72706 36706 72718
rect 47070 72770 47122 72782
rect 57138 72718 57150 72770
rect 57202 72718 57214 72770
rect 59602 72718 59614 72770
rect 59666 72767 59678 72770
rect 60162 72767 60174 72770
rect 59666 72721 60174 72767
rect 59666 72718 59678 72721
rect 60162 72718 60174 72721
rect 60226 72718 60238 72770
rect 47070 72706 47122 72718
rect 30942 72658 30994 72670
rect 30942 72594 30994 72606
rect 32622 72658 32674 72670
rect 32622 72594 32674 72606
rect 33070 72658 33122 72670
rect 33070 72594 33122 72606
rect 33406 72658 33458 72670
rect 33406 72594 33458 72606
rect 33854 72658 33906 72670
rect 43934 72658 43986 72670
rect 43138 72606 43150 72658
rect 43202 72606 43214 72658
rect 33854 72594 33906 72606
rect 43934 72594 43986 72606
rect 47182 72658 47234 72670
rect 55806 72658 55858 72670
rect 59390 72658 59442 72670
rect 52434 72606 52446 72658
rect 52498 72606 52510 72658
rect 54338 72606 54350 72658
rect 54402 72606 54414 72658
rect 56578 72606 56590 72658
rect 56642 72606 56654 72658
rect 47182 72594 47234 72606
rect 55806 72594 55858 72606
rect 59390 72594 59442 72606
rect 59838 72658 59890 72670
rect 59838 72594 59890 72606
rect 60286 72658 60338 72670
rect 60286 72594 60338 72606
rect 61294 72658 61346 72670
rect 61294 72594 61346 72606
rect 35086 72546 35138 72558
rect 35086 72482 35138 72494
rect 37774 72546 37826 72558
rect 41582 72546 41634 72558
rect 44046 72546 44098 72558
rect 39106 72494 39118 72546
rect 39170 72494 39182 72546
rect 40114 72494 40126 72546
rect 40178 72494 40190 72546
rect 42690 72494 42702 72546
rect 42754 72494 42766 72546
rect 37774 72482 37826 72494
rect 41582 72482 41634 72494
rect 44046 72482 44098 72494
rect 44494 72546 44546 72558
rect 44494 72482 44546 72494
rect 45614 72546 45666 72558
rect 49870 72546 49922 72558
rect 46162 72494 46174 72546
rect 46226 72494 46238 72546
rect 45614 72482 45666 72494
rect 49870 72482 49922 72494
rect 50094 72546 50146 72558
rect 52670 72546 52722 72558
rect 50418 72494 50430 72546
rect 50482 72494 50494 72546
rect 52098 72494 52110 72546
rect 52162 72494 52174 72546
rect 50094 72482 50146 72494
rect 52670 72482 52722 72494
rect 53454 72546 53506 72558
rect 55358 72546 55410 72558
rect 57822 72546 57874 72558
rect 59278 72546 59330 72558
rect 53890 72494 53902 72546
rect 53954 72494 53966 72546
rect 57026 72494 57038 72546
rect 57090 72494 57102 72546
rect 57474 72494 57486 72546
rect 57538 72494 57550 72546
rect 58034 72494 58046 72546
rect 58098 72494 58110 72546
rect 53454 72482 53506 72494
rect 55358 72482 55410 72494
rect 57822 72482 57874 72494
rect 59278 72482 59330 72494
rect 34414 72434 34466 72446
rect 34414 72370 34466 72382
rect 34526 72434 34578 72446
rect 34526 72370 34578 72382
rect 35198 72434 35250 72446
rect 35198 72370 35250 72382
rect 35982 72434 36034 72446
rect 35982 72370 36034 72382
rect 36542 72434 36594 72446
rect 36542 72370 36594 72382
rect 36654 72434 36706 72446
rect 36654 72370 36706 72382
rect 37438 72434 37490 72446
rect 41694 72434 41746 72446
rect 38882 72382 38894 72434
rect 38946 72382 38958 72434
rect 37438 72370 37490 72382
rect 41694 72370 41746 72382
rect 42254 72434 42306 72446
rect 42254 72370 42306 72382
rect 45502 72434 45554 72446
rect 45502 72370 45554 72382
rect 47742 72434 47794 72446
rect 47742 72370 47794 72382
rect 48414 72434 48466 72446
rect 48414 72370 48466 72382
rect 49310 72434 49362 72446
rect 49310 72370 49362 72382
rect 55022 72434 55074 72446
rect 55022 72370 55074 72382
rect 31950 72322 32002 72334
rect 31950 72258 32002 72270
rect 37662 72322 37714 72334
rect 41470 72322 41522 72334
rect 40226 72270 40238 72322
rect 40290 72270 40302 72322
rect 37662 72258 37714 72270
rect 41470 72258 41522 72270
rect 43822 72322 43874 72334
rect 43822 72258 43874 72270
rect 49982 72322 50034 72334
rect 49982 72258 50034 72270
rect 50878 72322 50930 72334
rect 50878 72258 50930 72270
rect 1344 72154 78624 72188
rect 1344 72102 19838 72154
rect 19890 72102 19942 72154
rect 19994 72102 20046 72154
rect 20098 72102 50558 72154
rect 50610 72102 50662 72154
rect 50714 72102 50766 72154
rect 50818 72102 78624 72154
rect 1344 72068 78624 72102
rect 33966 71986 34018 71998
rect 33966 71922 34018 71934
rect 34302 71986 34354 71998
rect 34302 71922 34354 71934
rect 35422 71986 35474 71998
rect 35422 71922 35474 71934
rect 36094 71986 36146 71998
rect 36094 71922 36146 71934
rect 36430 71986 36482 71998
rect 36430 71922 36482 71934
rect 37102 71986 37154 71998
rect 37102 71922 37154 71934
rect 37998 71986 38050 71998
rect 37998 71922 38050 71934
rect 41470 71986 41522 71998
rect 44942 71986 44994 71998
rect 43586 71934 43598 71986
rect 43650 71934 43662 71986
rect 41470 71922 41522 71934
rect 44942 71922 44994 71934
rect 45166 71986 45218 71998
rect 45166 71922 45218 71934
rect 45950 71986 46002 71998
rect 45950 71922 46002 71934
rect 46622 71986 46674 71998
rect 46622 71922 46674 71934
rect 47294 71986 47346 71998
rect 47294 71922 47346 71934
rect 47742 71986 47794 71998
rect 47742 71922 47794 71934
rect 48638 71986 48690 71998
rect 59054 71986 59106 71998
rect 53890 71934 53902 71986
rect 53954 71934 53966 71986
rect 56578 71934 56590 71986
rect 56642 71934 56654 71986
rect 48638 71922 48690 71934
rect 59054 71922 59106 71934
rect 59614 71986 59666 71998
rect 59614 71922 59666 71934
rect 34750 71874 34802 71886
rect 34750 71810 34802 71822
rect 36990 71874 37042 71886
rect 46062 71874 46114 71886
rect 52446 71874 52498 71886
rect 43474 71822 43486 71874
rect 43538 71822 43550 71874
rect 44146 71822 44158 71874
rect 44210 71822 44222 71874
rect 49746 71822 49758 71874
rect 49810 71822 49822 71874
rect 36990 71810 37042 71822
rect 46062 71810 46114 71822
rect 52446 71810 52498 71822
rect 52782 71874 52834 71886
rect 52782 71810 52834 71822
rect 55470 71874 55522 71886
rect 55470 71810 55522 71822
rect 58606 71874 58658 71886
rect 58606 71810 58658 71822
rect 45278 71762 45330 71774
rect 37762 71710 37774 71762
rect 37826 71710 37838 71762
rect 38770 71710 38782 71762
rect 38834 71710 38846 71762
rect 39106 71710 39118 71762
rect 39170 71710 39182 71762
rect 40450 71710 40462 71762
rect 40514 71710 40526 71762
rect 42130 71710 42142 71762
rect 42194 71710 42206 71762
rect 43026 71710 43038 71762
rect 43090 71710 43102 71762
rect 43810 71710 43822 71762
rect 43874 71710 43886 71762
rect 45278 71698 45330 71710
rect 45726 71762 45778 71774
rect 52558 71762 52610 71774
rect 50306 71710 50318 71762
rect 50370 71710 50382 71762
rect 51314 71710 51326 71762
rect 51378 71710 51390 71762
rect 45726 71698 45778 71710
rect 52558 71698 52610 71710
rect 52894 71762 52946 71774
rect 52894 71698 52946 71710
rect 54238 71762 54290 71774
rect 54238 71698 54290 71710
rect 54462 71762 54514 71774
rect 56030 71762 56082 71774
rect 55234 71710 55246 71762
rect 55298 71710 55310 71762
rect 58034 71710 58046 71762
rect 58098 71710 58110 71762
rect 54462 71698 54514 71710
rect 56030 71698 56082 71710
rect 48190 71650 48242 71662
rect 39218 71598 39230 71650
rect 39282 71598 39294 71650
rect 40338 71598 40350 71650
rect 40402 71598 40414 71650
rect 51762 71598 51774 71650
rect 51826 71598 51838 71650
rect 57810 71598 57822 71650
rect 57874 71598 57886 71650
rect 48190 71586 48242 71598
rect 56254 71538 56306 71550
rect 40226 71486 40238 71538
rect 40290 71486 40302 71538
rect 48178 71486 48190 71538
rect 48242 71535 48254 71538
rect 48626 71535 48638 71538
rect 48242 71489 48638 71535
rect 48242 71486 48254 71489
rect 48626 71486 48638 71489
rect 48690 71486 48702 71538
rect 56254 71474 56306 71486
rect 1344 71370 78624 71404
rect 1344 71318 4478 71370
rect 4530 71318 4582 71370
rect 4634 71318 4686 71370
rect 4738 71318 35198 71370
rect 35250 71318 35302 71370
rect 35354 71318 35406 71370
rect 35458 71318 65918 71370
rect 65970 71318 66022 71370
rect 66074 71318 66126 71370
rect 66178 71318 78624 71370
rect 1344 71284 78624 71318
rect 39678 71202 39730 71214
rect 33618 71150 33630 71202
rect 33682 71199 33694 71202
rect 34738 71199 34750 71202
rect 33682 71153 34750 71199
rect 33682 71150 33694 71153
rect 34738 71150 34750 71153
rect 34802 71150 34814 71202
rect 39106 71150 39118 71202
rect 39170 71150 39182 71202
rect 39678 71138 39730 71150
rect 40014 71202 40066 71214
rect 49186 71150 49198 71202
rect 49250 71199 49262 71202
rect 50306 71199 50318 71202
rect 49250 71153 50318 71199
rect 49250 71150 49262 71153
rect 50306 71150 50318 71153
rect 50370 71150 50382 71202
rect 54450 71150 54462 71202
rect 54514 71199 54526 71202
rect 54674 71199 54686 71202
rect 54514 71153 54686 71199
rect 54514 71150 54526 71153
rect 54674 71150 54686 71153
rect 54738 71199 54750 71202
rect 55010 71199 55022 71202
rect 54738 71153 55022 71199
rect 54738 71150 54750 71153
rect 55010 71150 55022 71153
rect 55074 71199 55086 71202
rect 55234 71199 55246 71202
rect 55074 71153 55246 71199
rect 55074 71150 55086 71153
rect 55234 71150 55246 71153
rect 55298 71150 55310 71202
rect 40014 71138 40066 71150
rect 34750 71090 34802 71102
rect 34750 71026 34802 71038
rect 35310 71090 35362 71102
rect 35310 71026 35362 71038
rect 36430 71090 36482 71102
rect 36430 71026 36482 71038
rect 36878 71090 36930 71102
rect 36878 71026 36930 71038
rect 37662 71090 37714 71102
rect 37662 71026 37714 71038
rect 38558 71090 38610 71102
rect 45390 71090 45442 71102
rect 41010 71038 41022 71090
rect 41074 71038 41086 71090
rect 42354 71038 42366 71090
rect 42418 71038 42430 71090
rect 44146 71038 44158 71090
rect 44210 71038 44222 71090
rect 38558 71026 38610 71038
rect 45390 71026 45442 71038
rect 45950 71090 46002 71102
rect 45950 71026 46002 71038
rect 46734 71090 46786 71102
rect 46734 71026 46786 71038
rect 47406 71090 47458 71102
rect 47406 71026 47458 71038
rect 47854 71090 47906 71102
rect 47854 71026 47906 71038
rect 48302 71090 48354 71102
rect 48302 71026 48354 71038
rect 49198 71090 49250 71102
rect 49198 71026 49250 71038
rect 49758 71090 49810 71102
rect 49758 71026 49810 71038
rect 50318 71090 50370 71102
rect 50318 71026 50370 71038
rect 50878 71090 50930 71102
rect 50878 71026 50930 71038
rect 54686 71090 54738 71102
rect 54686 71026 54738 71038
rect 55246 71090 55298 71102
rect 55246 71026 55298 71038
rect 55694 71090 55746 71102
rect 55694 71026 55746 71038
rect 58942 71090 58994 71102
rect 58942 71026 58994 71038
rect 38782 70978 38834 70990
rect 41806 70978 41858 70990
rect 48750 70978 48802 70990
rect 39666 70926 39678 70978
rect 39730 70926 39742 70978
rect 41234 70926 41246 70978
rect 41298 70926 41310 70978
rect 42802 70926 42814 70978
rect 42866 70926 42878 70978
rect 44482 70926 44494 70978
rect 44546 70926 44558 70978
rect 57026 70926 57038 70978
rect 57090 70926 57102 70978
rect 38782 70914 38834 70926
rect 41806 70914 41858 70926
rect 48750 70914 48802 70926
rect 38110 70866 38162 70878
rect 38110 70802 38162 70814
rect 51550 70866 51602 70878
rect 51550 70802 51602 70814
rect 52222 70866 52274 70878
rect 52222 70802 52274 70814
rect 53566 70866 53618 70878
rect 56914 70814 56926 70866
rect 56978 70814 56990 70866
rect 58258 70814 58270 70866
rect 58322 70814 58334 70866
rect 53566 70802 53618 70814
rect 46286 70754 46338 70766
rect 46286 70690 46338 70702
rect 54126 70754 54178 70766
rect 58146 70702 58158 70754
rect 58210 70702 58222 70754
rect 54126 70690 54178 70702
rect 1344 70586 78624 70620
rect 1344 70534 19838 70586
rect 19890 70534 19942 70586
rect 19994 70534 20046 70586
rect 20098 70534 50558 70586
rect 50610 70534 50662 70586
rect 50714 70534 50766 70586
rect 50818 70534 78624 70586
rect 1344 70500 78624 70534
rect 37102 70418 37154 70430
rect 37102 70354 37154 70366
rect 37998 70418 38050 70430
rect 37998 70354 38050 70366
rect 39006 70418 39058 70430
rect 39006 70354 39058 70366
rect 39566 70418 39618 70430
rect 39566 70354 39618 70366
rect 41582 70418 41634 70430
rect 41582 70354 41634 70366
rect 42702 70418 42754 70430
rect 44718 70418 44770 70430
rect 43586 70366 43598 70418
rect 43650 70366 43662 70418
rect 42702 70354 42754 70366
rect 44718 70354 44770 70366
rect 45054 70418 45106 70430
rect 45054 70354 45106 70366
rect 45502 70418 45554 70430
rect 45502 70354 45554 70366
rect 46398 70418 46450 70430
rect 46398 70354 46450 70366
rect 46846 70418 46898 70430
rect 46846 70354 46898 70366
rect 47182 70418 47234 70430
rect 47182 70354 47234 70366
rect 48414 70418 48466 70430
rect 48414 70354 48466 70366
rect 50430 70418 50482 70430
rect 50430 70354 50482 70366
rect 51326 70418 51378 70430
rect 51326 70354 51378 70366
rect 51774 70418 51826 70430
rect 51774 70354 51826 70366
rect 52222 70418 52274 70430
rect 52222 70354 52274 70366
rect 52670 70418 52722 70430
rect 52670 70354 52722 70366
rect 53118 70418 53170 70430
rect 53118 70354 53170 70366
rect 53566 70418 53618 70430
rect 53566 70354 53618 70366
rect 54574 70418 54626 70430
rect 54574 70354 54626 70366
rect 55022 70418 55074 70430
rect 55570 70366 55582 70418
rect 55634 70415 55646 70418
rect 56354 70415 56366 70418
rect 55634 70369 56366 70415
rect 55634 70366 55646 70369
rect 56354 70366 56366 70369
rect 56418 70366 56430 70418
rect 55022 70354 55074 70366
rect 37438 70306 37490 70318
rect 37438 70242 37490 70254
rect 39678 70306 39730 70318
rect 39678 70242 39730 70254
rect 40350 70306 40402 70318
rect 40350 70242 40402 70254
rect 40798 70306 40850 70318
rect 40798 70242 40850 70254
rect 43038 70306 43090 70318
rect 43038 70242 43090 70254
rect 55470 70306 55522 70318
rect 55470 70242 55522 70254
rect 40238 70194 40290 70206
rect 40238 70130 40290 70142
rect 42366 70194 42418 70206
rect 42366 70130 42418 70142
rect 42814 70194 42866 70206
rect 42814 70130 42866 70142
rect 43934 70194 43986 70206
rect 43934 70130 43986 70142
rect 44158 70194 44210 70206
rect 44158 70130 44210 70142
rect 38334 70082 38386 70094
rect 38334 70018 38386 70030
rect 37538 69918 37550 69970
rect 37602 69967 37614 69970
rect 38322 69967 38334 69970
rect 37602 69921 38334 69967
rect 37602 69918 37614 69921
rect 38322 69918 38334 69921
rect 38386 69918 38398 69970
rect 1344 69802 78624 69836
rect 1344 69750 4478 69802
rect 4530 69750 4582 69802
rect 4634 69750 4686 69802
rect 4738 69750 35198 69802
rect 35250 69750 35302 69802
rect 35354 69750 35406 69802
rect 35458 69750 65918 69802
rect 65970 69750 66022 69802
rect 66074 69750 66126 69802
rect 66178 69750 78624 69802
rect 1344 69716 78624 69750
rect 38322 69582 38334 69634
rect 38386 69631 38398 69634
rect 39778 69631 39790 69634
rect 38386 69585 39790 69631
rect 38386 69582 38398 69585
rect 39778 69582 39790 69585
rect 39842 69582 39854 69634
rect 39790 69522 39842 69534
rect 39790 69458 39842 69470
rect 40350 69522 40402 69534
rect 40350 69458 40402 69470
rect 40798 69522 40850 69534
rect 40798 69458 40850 69470
rect 46174 69522 46226 69534
rect 46174 69458 46226 69470
rect 46622 69522 46674 69534
rect 46622 69458 46674 69470
rect 52334 69522 52386 69534
rect 52334 69458 52386 69470
rect 52782 69522 52834 69534
rect 52782 69458 52834 69470
rect 1344 69018 78624 69052
rect 1344 68966 19838 69018
rect 19890 68966 19942 69018
rect 19994 68966 20046 69018
rect 20098 68966 50558 69018
rect 50610 68966 50662 69018
rect 50714 68966 50766 69018
rect 50818 68966 78624 69018
rect 1344 68932 78624 68966
rect 1344 68234 78624 68268
rect 1344 68182 4478 68234
rect 4530 68182 4582 68234
rect 4634 68182 4686 68234
rect 4738 68182 35198 68234
rect 35250 68182 35302 68234
rect 35354 68182 35406 68234
rect 35458 68182 65918 68234
rect 65970 68182 66022 68234
rect 66074 68182 66126 68234
rect 66178 68182 78624 68234
rect 1344 68148 78624 68182
rect 1344 67450 78624 67484
rect 1344 67398 19838 67450
rect 19890 67398 19942 67450
rect 19994 67398 20046 67450
rect 20098 67398 50558 67450
rect 50610 67398 50662 67450
rect 50714 67398 50766 67450
rect 50818 67398 78624 67450
rect 1344 67364 78624 67398
rect 1344 66666 78624 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 35198 66666
rect 35250 66614 35302 66666
rect 35354 66614 35406 66666
rect 35458 66614 65918 66666
rect 65970 66614 66022 66666
rect 66074 66614 66126 66666
rect 66178 66614 78624 66666
rect 1344 66580 78624 66614
rect 1344 65882 78624 65916
rect 1344 65830 19838 65882
rect 19890 65830 19942 65882
rect 19994 65830 20046 65882
rect 20098 65830 50558 65882
rect 50610 65830 50662 65882
rect 50714 65830 50766 65882
rect 50818 65830 78624 65882
rect 1344 65796 78624 65830
rect 1344 65098 78624 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 35198 65098
rect 35250 65046 35302 65098
rect 35354 65046 35406 65098
rect 35458 65046 65918 65098
rect 65970 65046 66022 65098
rect 66074 65046 66126 65098
rect 66178 65046 78624 65098
rect 1344 65012 78624 65046
rect 1344 64314 78624 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 50558 64314
rect 50610 64262 50662 64314
rect 50714 64262 50766 64314
rect 50818 64262 78624 64314
rect 1344 64228 78624 64262
rect 1344 63530 78624 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 65918 63530
rect 65970 63478 66022 63530
rect 66074 63478 66126 63530
rect 66178 63478 78624 63530
rect 1344 63444 78624 63478
rect 1344 62746 78624 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 50558 62746
rect 50610 62694 50662 62746
rect 50714 62694 50766 62746
rect 50818 62694 78624 62746
rect 1344 62660 78624 62694
rect 1344 61962 78624 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 65918 61962
rect 65970 61910 66022 61962
rect 66074 61910 66126 61962
rect 66178 61910 78624 61962
rect 1344 61876 78624 61910
rect 1344 61178 78624 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 50558 61178
rect 50610 61126 50662 61178
rect 50714 61126 50766 61178
rect 50818 61126 78624 61178
rect 1344 61092 78624 61126
rect 1344 60394 78624 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 65918 60394
rect 65970 60342 66022 60394
rect 66074 60342 66126 60394
rect 66178 60342 78624 60394
rect 1344 60308 78624 60342
rect 1344 59610 78624 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 50558 59610
rect 50610 59558 50662 59610
rect 50714 59558 50766 59610
rect 50818 59558 78624 59610
rect 1344 59524 78624 59558
rect 1344 58826 78624 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 65918 58826
rect 65970 58774 66022 58826
rect 66074 58774 66126 58826
rect 66178 58774 78624 58826
rect 1344 58740 78624 58774
rect 1344 58042 78624 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 50558 58042
rect 50610 57990 50662 58042
rect 50714 57990 50766 58042
rect 50818 57990 78624 58042
rect 1344 57956 78624 57990
rect 1344 57258 78624 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 65918 57258
rect 65970 57206 66022 57258
rect 66074 57206 66126 57258
rect 66178 57206 78624 57258
rect 1344 57172 78624 57206
rect 1344 56474 78624 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 78624 56474
rect 1344 56388 78624 56422
rect 1344 55690 78624 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 65918 55690
rect 65970 55638 66022 55690
rect 66074 55638 66126 55690
rect 66178 55638 78624 55690
rect 1344 55604 78624 55638
rect 1344 54906 78624 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 78624 54906
rect 1344 54820 78624 54854
rect 1344 54122 78624 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 65918 54122
rect 65970 54070 66022 54122
rect 66074 54070 66126 54122
rect 66178 54070 78624 54122
rect 1344 54036 78624 54070
rect 1344 53338 78624 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 78624 53338
rect 1344 53252 78624 53286
rect 1344 52554 78624 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 65918 52554
rect 65970 52502 66022 52554
rect 66074 52502 66126 52554
rect 66178 52502 78624 52554
rect 1344 52468 78624 52502
rect 1344 51770 78624 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 78624 51770
rect 1344 51684 78624 51718
rect 1344 50986 78624 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 65918 50986
rect 65970 50934 66022 50986
rect 66074 50934 66126 50986
rect 66178 50934 78624 50986
rect 1344 50900 78624 50934
rect 1344 50202 78624 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 78624 50202
rect 1344 50116 78624 50150
rect 1344 49418 78624 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 65918 49418
rect 65970 49366 66022 49418
rect 66074 49366 66126 49418
rect 66178 49366 78624 49418
rect 1344 49332 78624 49366
rect 1344 48634 78624 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 78624 48634
rect 1344 48548 78624 48582
rect 1344 47850 78624 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 65918 47850
rect 65970 47798 66022 47850
rect 66074 47798 66126 47850
rect 66178 47798 78624 47850
rect 1344 47764 78624 47798
rect 1344 47066 78624 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 78624 47066
rect 1344 46980 78624 47014
rect 1344 46282 78624 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 65918 46282
rect 65970 46230 66022 46282
rect 66074 46230 66126 46282
rect 66178 46230 78624 46282
rect 1344 46196 78624 46230
rect 1344 45498 78624 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 78624 45498
rect 1344 45412 78624 45446
rect 1344 44714 78624 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 65918 44714
rect 65970 44662 66022 44714
rect 66074 44662 66126 44714
rect 66178 44662 78624 44714
rect 1344 44628 78624 44662
rect 1344 43930 78624 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 78624 43930
rect 1344 43844 78624 43878
rect 1344 43146 78624 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 65918 43146
rect 65970 43094 66022 43146
rect 66074 43094 66126 43146
rect 66178 43094 78624 43146
rect 1344 43060 78624 43094
rect 1344 42362 78624 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 78624 42362
rect 1344 42276 78624 42310
rect 1344 41578 78624 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 65918 41578
rect 65970 41526 66022 41578
rect 66074 41526 66126 41578
rect 66178 41526 78624 41578
rect 1344 41492 78624 41526
rect 1344 40794 78624 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 78624 40794
rect 1344 40708 78624 40742
rect 1344 40010 78624 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 65918 40010
rect 65970 39958 66022 40010
rect 66074 39958 66126 40010
rect 66178 39958 78624 40010
rect 1344 39924 78624 39958
rect 1344 39226 78624 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 78624 39226
rect 1344 39140 78624 39174
rect 1344 38442 78624 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 65918 38442
rect 65970 38390 66022 38442
rect 66074 38390 66126 38442
rect 66178 38390 78624 38442
rect 1344 38356 78624 38390
rect 1344 37658 78624 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 78624 37658
rect 1344 37572 78624 37606
rect 1344 36874 78624 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 65918 36874
rect 65970 36822 66022 36874
rect 66074 36822 66126 36874
rect 66178 36822 78624 36874
rect 1344 36788 78624 36822
rect 1344 36090 78624 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 78624 36090
rect 1344 36004 78624 36038
rect 1344 35306 78624 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 65918 35306
rect 65970 35254 66022 35306
rect 66074 35254 66126 35306
rect 66178 35254 78624 35306
rect 1344 35220 78624 35254
rect 1344 34522 78624 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 78624 34522
rect 1344 34436 78624 34470
rect 1344 33738 78624 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 65918 33738
rect 65970 33686 66022 33738
rect 66074 33686 66126 33738
rect 66178 33686 78624 33738
rect 1344 33652 78624 33686
rect 1344 32954 78624 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 78624 32954
rect 1344 32868 78624 32902
rect 1344 32170 78624 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 65918 32170
rect 65970 32118 66022 32170
rect 66074 32118 66126 32170
rect 66178 32118 78624 32170
rect 1344 32084 78624 32118
rect 1344 31386 78624 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 78624 31386
rect 1344 31300 78624 31334
rect 1344 30602 78624 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 65918 30602
rect 65970 30550 66022 30602
rect 66074 30550 66126 30602
rect 66178 30550 78624 30602
rect 1344 30516 78624 30550
rect 1344 29818 78624 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 78624 29818
rect 1344 29732 78624 29766
rect 1344 29034 78624 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 65918 29034
rect 65970 28982 66022 29034
rect 66074 28982 66126 29034
rect 66178 28982 78624 29034
rect 1344 28948 78624 28982
rect 1344 28250 78624 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 78624 28250
rect 1344 28164 78624 28198
rect 1344 27466 78624 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 65918 27466
rect 65970 27414 66022 27466
rect 66074 27414 66126 27466
rect 66178 27414 78624 27466
rect 1344 27380 78624 27414
rect 1344 26682 78624 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 78624 26682
rect 1344 26596 78624 26630
rect 1344 25898 78624 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 65918 25898
rect 65970 25846 66022 25898
rect 66074 25846 66126 25898
rect 66178 25846 78624 25898
rect 1344 25812 78624 25846
rect 1344 25114 78624 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 78624 25114
rect 1344 25028 78624 25062
rect 1344 24330 78624 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 65918 24330
rect 65970 24278 66022 24330
rect 66074 24278 66126 24330
rect 66178 24278 78624 24330
rect 1344 24244 78624 24278
rect 1344 23546 78624 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 78624 23546
rect 1344 23460 78624 23494
rect 1344 22762 78624 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 65918 22762
rect 65970 22710 66022 22762
rect 66074 22710 66126 22762
rect 66178 22710 78624 22762
rect 1344 22676 78624 22710
rect 1344 21978 78624 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 78624 21978
rect 1344 21892 78624 21926
rect 1344 21194 78624 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 65918 21194
rect 65970 21142 66022 21194
rect 66074 21142 66126 21194
rect 66178 21142 78624 21194
rect 1344 21108 78624 21142
rect 1344 20410 78624 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 78624 20410
rect 1344 20324 78624 20358
rect 1344 19626 78624 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 65918 19626
rect 65970 19574 66022 19626
rect 66074 19574 66126 19626
rect 66178 19574 78624 19626
rect 1344 19540 78624 19574
rect 1344 18842 78624 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 78624 18842
rect 1344 18756 78624 18790
rect 1344 18058 78624 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 65918 18058
rect 65970 18006 66022 18058
rect 66074 18006 66126 18058
rect 66178 18006 78624 18058
rect 1344 17972 78624 18006
rect 1344 17274 78624 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 78624 17274
rect 1344 17188 78624 17222
rect 1344 16490 78624 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 65918 16490
rect 65970 16438 66022 16490
rect 66074 16438 66126 16490
rect 66178 16438 78624 16490
rect 1344 16404 78624 16438
rect 1344 15706 78624 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 78624 15706
rect 1344 15620 78624 15654
rect 1344 14922 78624 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 65918 14922
rect 65970 14870 66022 14922
rect 66074 14870 66126 14922
rect 66178 14870 78624 14922
rect 1344 14836 78624 14870
rect 1344 14138 78624 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 78624 14138
rect 1344 14052 78624 14086
rect 1344 13354 78624 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 65918 13354
rect 65970 13302 66022 13354
rect 66074 13302 66126 13354
rect 66178 13302 78624 13354
rect 1344 13268 78624 13302
rect 1344 12570 78624 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 78624 12570
rect 1344 12484 78624 12518
rect 1344 11786 78624 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 65918 11786
rect 65970 11734 66022 11786
rect 66074 11734 66126 11786
rect 66178 11734 78624 11786
rect 1344 11700 78624 11734
rect 1344 11002 78624 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 78624 11002
rect 1344 10916 78624 10950
rect 1344 10218 78624 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 65918 10218
rect 65970 10166 66022 10218
rect 66074 10166 66126 10218
rect 66178 10166 78624 10218
rect 1344 10132 78624 10166
rect 1344 9434 78624 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 78624 9434
rect 1344 9348 78624 9382
rect 1344 8650 78624 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 65918 8650
rect 65970 8598 66022 8650
rect 66074 8598 66126 8650
rect 66178 8598 78624 8650
rect 1344 8564 78624 8598
rect 1344 7866 78624 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 78624 7866
rect 1344 7780 78624 7814
rect 1344 7082 78624 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 65918 7082
rect 65970 7030 66022 7082
rect 66074 7030 66126 7082
rect 66178 7030 78624 7082
rect 1344 6996 78624 7030
rect 1344 6298 78624 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 78624 6298
rect 1344 6212 78624 6246
rect 1344 5514 78624 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 65918 5514
rect 65970 5462 66022 5514
rect 66074 5462 66126 5514
rect 66178 5462 78624 5514
rect 1344 5428 78624 5462
rect 1344 4730 78624 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 78624 4730
rect 1344 4644 78624 4678
rect 13918 4450 13970 4462
rect 13918 4386 13970 4398
rect 17950 4450 18002 4462
rect 17950 4386 18002 4398
rect 24670 4450 24722 4462
rect 24670 4386 24722 4398
rect 29374 4450 29426 4462
rect 29374 4386 29426 4398
rect 32510 4450 32562 4462
rect 32510 4386 32562 4398
rect 37214 4450 37266 4462
rect 37214 4386 37266 4398
rect 51326 4450 51378 4462
rect 51326 4386 51378 4398
rect 55358 4450 55410 4462
rect 55358 4386 55410 4398
rect 59390 4450 59442 4462
rect 59390 4386 59442 4398
rect 63422 4450 63474 4462
rect 63422 4386 63474 4398
rect 70814 4450 70866 4462
rect 70814 4386 70866 4398
rect 73390 4450 73442 4462
rect 73390 4386 73442 4398
rect 74062 4450 74114 4462
rect 74062 4386 74114 4398
rect 1344 3946 78624 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 65918 3946
rect 65970 3894 66022 3946
rect 66074 3894 66126 3946
rect 66178 3894 78624 3946
rect 1344 3860 78624 3894
rect 6974 3330 7026 3342
rect 6974 3266 7026 3278
rect 8094 3330 8146 3342
rect 8094 3266 8146 3278
rect 8878 3330 8930 3342
rect 8878 3266 8930 3278
rect 9998 3330 10050 3342
rect 9998 3266 10050 3278
rect 10782 3330 10834 3342
rect 10782 3266 10834 3278
rect 11454 3330 11506 3342
rect 11454 3266 11506 3278
rect 12126 3330 12178 3342
rect 12126 3266 12178 3278
rect 12798 3330 12850 3342
rect 12798 3266 12850 3278
rect 14030 3330 14082 3342
rect 14030 3266 14082 3278
rect 14702 3330 14754 3342
rect 14702 3266 14754 3278
rect 15374 3330 15426 3342
rect 15374 3266 15426 3278
rect 16046 3330 16098 3342
rect 16046 3266 16098 3278
rect 16718 3330 16770 3342
rect 16718 3266 16770 3278
rect 17950 3330 18002 3342
rect 17950 3266 18002 3278
rect 18622 3330 18674 3342
rect 18622 3266 18674 3278
rect 19294 3330 19346 3342
rect 19294 3266 19346 3278
rect 19966 3330 20018 3342
rect 19966 3266 20018 3278
rect 20638 3330 20690 3342
rect 20638 3266 20690 3278
rect 21758 3330 21810 3342
rect 21758 3266 21810 3278
rect 22430 3330 22482 3342
rect 22430 3266 22482 3278
rect 23102 3330 23154 3342
rect 23102 3266 23154 3278
rect 23774 3330 23826 3342
rect 23774 3266 23826 3278
rect 24558 3330 24610 3342
rect 24558 3266 24610 3278
rect 25790 3330 25842 3342
rect 25790 3266 25842 3278
rect 26462 3330 26514 3342
rect 26462 3266 26514 3278
rect 27134 3330 27186 3342
rect 27134 3266 27186 3278
rect 27806 3330 27858 3342
rect 27806 3266 27858 3278
rect 28478 3330 28530 3342
rect 28478 3266 28530 3278
rect 29710 3330 29762 3342
rect 29710 3266 29762 3278
rect 30270 3330 30322 3342
rect 30270 3266 30322 3278
rect 30942 3330 30994 3342
rect 30942 3266 30994 3278
rect 31614 3330 31666 3342
rect 31614 3266 31666 3278
rect 32398 3330 32450 3342
rect 32398 3266 32450 3278
rect 33630 3330 33682 3342
rect 33630 3266 33682 3278
rect 34302 3330 34354 3342
rect 34302 3266 34354 3278
rect 34974 3330 35026 3342
rect 34974 3266 35026 3278
rect 35646 3330 35698 3342
rect 35646 3266 35698 3278
rect 36318 3330 36370 3342
rect 36318 3266 36370 3278
rect 37550 3330 37602 3342
rect 37550 3266 37602 3278
rect 38222 3330 38274 3342
rect 38222 3266 38274 3278
rect 38894 3330 38946 3342
rect 38894 3266 38946 3278
rect 39566 3330 39618 3342
rect 39566 3266 39618 3278
rect 40238 3330 40290 3342
rect 40238 3266 40290 3278
rect 41246 3330 41298 3342
rect 41246 3266 41298 3278
rect 41918 3330 41970 3342
rect 41918 3266 41970 3278
rect 42590 3330 42642 3342
rect 42590 3266 42642 3278
rect 43262 3330 43314 3342
rect 43262 3266 43314 3278
rect 43934 3330 43986 3342
rect 43934 3266 43986 3278
rect 44942 3330 44994 3342
rect 44942 3266 44994 3278
rect 45614 3330 45666 3342
rect 45614 3266 45666 3278
rect 46286 3330 46338 3342
rect 46286 3266 46338 3278
rect 46958 3330 47010 3342
rect 46958 3266 47010 3278
rect 47630 3330 47682 3342
rect 47630 3266 47682 3278
rect 48862 3330 48914 3342
rect 48862 3266 48914 3278
rect 49534 3330 49586 3342
rect 49534 3266 49586 3278
rect 50206 3330 50258 3342
rect 50206 3266 50258 3278
rect 50878 3330 50930 3342
rect 50878 3266 50930 3278
rect 51550 3330 51602 3342
rect 51550 3266 51602 3278
rect 52782 3330 52834 3342
rect 52782 3266 52834 3278
rect 53454 3330 53506 3342
rect 53454 3266 53506 3278
rect 54126 3330 54178 3342
rect 54126 3266 54178 3278
rect 54798 3330 54850 3342
rect 54798 3266 54850 3278
rect 55470 3330 55522 3342
rect 55470 3266 55522 3278
rect 56702 3330 56754 3342
rect 56702 3266 56754 3278
rect 57374 3330 57426 3342
rect 57374 3266 57426 3278
rect 58046 3330 58098 3342
rect 58046 3266 58098 3278
rect 58718 3330 58770 3342
rect 58718 3266 58770 3278
rect 59390 3330 59442 3342
rect 59390 3266 59442 3278
rect 60622 3330 60674 3342
rect 60622 3266 60674 3278
rect 61294 3330 61346 3342
rect 61294 3266 61346 3278
rect 61966 3330 62018 3342
rect 61966 3266 62018 3278
rect 62638 3330 62690 3342
rect 62638 3266 62690 3278
rect 63310 3330 63362 3342
rect 63310 3266 63362 3278
rect 64542 3330 64594 3342
rect 64542 3266 64594 3278
rect 65214 3330 65266 3342
rect 65214 3266 65266 3278
rect 65886 3330 65938 3342
rect 65886 3266 65938 3278
rect 66558 3330 66610 3342
rect 66558 3266 66610 3278
rect 67230 3330 67282 3342
rect 67230 3266 67282 3278
rect 68462 3330 68514 3342
rect 68462 3266 68514 3278
rect 69134 3330 69186 3342
rect 69134 3266 69186 3278
rect 69806 3330 69858 3342
rect 69806 3266 69858 3278
rect 70478 3330 70530 3342
rect 70478 3266 70530 3278
rect 71150 3330 71202 3342
rect 71150 3266 71202 3278
rect 72382 3330 72434 3342
rect 72382 3266 72434 3278
rect 73054 3330 73106 3342
rect 73054 3266 73106 3278
rect 73726 3330 73778 3342
rect 73726 3266 73778 3278
rect 74398 3330 74450 3342
rect 74398 3266 74450 3278
rect 1344 3162 78624 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 78624 3162
rect 1344 3076 78624 3110
rect 46386 1822 46398 1874
rect 46450 1871 46462 1874
rect 46946 1871 46958 1874
rect 46450 1825 46958 1871
rect 46450 1822 46462 1825
rect 46946 1822 46958 1825
rect 47010 1822 47022 1874
rect 57810 1822 57822 1874
rect 57874 1871 57886 1874
rect 58706 1871 58718 1874
rect 57874 1825 58718 1871
rect 57874 1822 57886 1825
rect 58706 1822 58718 1825
rect 58770 1822 58782 1874
rect 61170 1822 61182 1874
rect 61234 1871 61246 1874
rect 61954 1871 61966 1874
rect 61234 1825 61966 1871
rect 61234 1822 61246 1825
rect 61954 1822 61966 1825
rect 62018 1822 62030 1874
rect 64642 1822 64654 1874
rect 64706 1871 64718 1874
rect 65202 1871 65214 1874
rect 64706 1825 65214 1871
rect 64706 1822 64718 1825
rect 65202 1822 65214 1825
rect 65266 1822 65278 1874
rect 65874 1822 65886 1874
rect 65938 1871 65950 1874
rect 66546 1871 66558 1874
rect 65938 1825 66558 1871
rect 65938 1822 65950 1825
rect 66546 1822 66558 1825
rect 66610 1822 66622 1874
rect 24546 1710 24558 1762
rect 24610 1759 24622 1762
rect 25106 1759 25118 1762
rect 24610 1713 25118 1759
rect 24610 1710 24622 1713
rect 25106 1710 25118 1713
rect 25170 1710 25182 1762
rect 32386 1710 32398 1762
rect 32450 1759 32462 1762
rect 32946 1759 32958 1762
rect 32450 1713 32958 1759
rect 32450 1710 32462 1713
rect 32946 1710 32958 1713
rect 33010 1710 33022 1762
rect 44370 1710 44382 1762
rect 44434 1759 44446 1762
rect 44930 1759 44942 1762
rect 44434 1713 44942 1759
rect 44434 1710 44446 1713
rect 44930 1710 44942 1713
rect 44994 1710 45006 1762
rect 45714 1710 45726 1762
rect 45778 1759 45790 1762
rect 46274 1759 46286 1762
rect 45778 1713 46286 1759
rect 45778 1710 45790 1713
rect 46274 1710 46286 1713
rect 46338 1710 46350 1762
rect 47058 1710 47070 1762
rect 47122 1759 47134 1762
rect 47618 1759 47630 1762
rect 47122 1713 47630 1759
rect 47122 1710 47134 1713
rect 47618 1710 47630 1713
rect 47682 1710 47694 1762
rect 49074 1710 49086 1762
rect 49138 1759 49150 1762
rect 50194 1759 50206 1762
rect 49138 1713 50206 1759
rect 49138 1710 49150 1713
rect 50194 1710 50206 1713
rect 50258 1710 50270 1762
rect 50418 1710 50430 1762
rect 50482 1759 50494 1762
rect 51538 1759 51550 1762
rect 50482 1713 51550 1759
rect 50482 1710 50494 1713
rect 51538 1710 51550 1713
rect 51602 1710 51614 1762
rect 52434 1710 52446 1762
rect 52498 1759 52510 1762
rect 53442 1759 53454 1762
rect 52498 1713 53454 1759
rect 52498 1710 52510 1713
rect 53442 1710 53454 1713
rect 53506 1710 53518 1762
rect 53778 1710 53790 1762
rect 53842 1759 53854 1762
rect 54786 1759 54798 1762
rect 53842 1713 54798 1759
rect 53842 1710 53854 1713
rect 54786 1710 54798 1713
rect 54850 1710 54862 1762
rect 55794 1710 55806 1762
rect 55858 1759 55870 1762
rect 56690 1759 56702 1762
rect 55858 1713 56702 1759
rect 55858 1710 55870 1713
rect 56690 1710 56702 1713
rect 56754 1710 56766 1762
rect 57138 1710 57150 1762
rect 57202 1759 57214 1762
rect 58034 1759 58046 1762
rect 57202 1713 58046 1759
rect 57202 1710 57214 1713
rect 58034 1710 58046 1713
rect 58098 1710 58110 1762
rect 60498 1710 60510 1762
rect 60562 1759 60574 1762
rect 61282 1759 61294 1762
rect 60562 1713 61294 1759
rect 60562 1710 60574 1713
rect 61282 1710 61294 1713
rect 61346 1710 61358 1762
rect 62514 1710 62526 1762
rect 62578 1759 62590 1762
rect 63298 1759 63310 1762
rect 62578 1713 63310 1759
rect 62578 1710 62590 1713
rect 63298 1710 63310 1713
rect 63362 1710 63374 1762
rect 63858 1710 63870 1762
rect 63922 1759 63934 1762
rect 64530 1759 64542 1762
rect 63922 1713 64542 1759
rect 63922 1710 63934 1713
rect 64530 1710 64542 1713
rect 64594 1710 64606 1762
rect 67218 1710 67230 1762
rect 67282 1759 67294 1762
rect 68450 1759 68462 1762
rect 67282 1713 68462 1759
rect 67282 1710 67294 1713
rect 68450 1710 68462 1713
rect 68514 1710 68526 1762
rect 69234 1710 69246 1762
rect 69298 1759 69310 1762
rect 70466 1759 70478 1762
rect 69298 1713 70478 1759
rect 69298 1710 69310 1713
rect 70466 1710 70478 1713
rect 70530 1710 70542 1762
rect 72594 1710 72606 1762
rect 72658 1759 72670 1762
rect 73714 1759 73726 1762
rect 72658 1713 73726 1759
rect 72658 1710 72670 1713
rect 73714 1710 73726 1713
rect 73778 1710 73790 1762
<< via1 >>
rect 74174 77198 74226 77250
rect 75294 77198 75346 77250
rect 32398 76974 32450 77026
rect 33294 76974 33346 77026
rect 37886 76974 37938 77026
rect 38782 76974 38834 77026
rect 45390 76974 45442 77026
rect 46734 76974 46786 77026
rect 48078 76974 48130 77026
rect 48638 76974 48690 77026
rect 60734 76974 60786 77026
rect 61294 76974 61346 77026
rect 76190 76974 76242 77026
rect 76974 76974 77026 77026
rect 19838 76806 19890 76858
rect 19942 76806 19994 76858
rect 20046 76806 20098 76858
rect 50558 76806 50610 76858
rect 50662 76806 50714 76858
rect 50766 76806 50818 76858
rect 3838 76638 3890 76690
rect 4958 76638 5010 76690
rect 7870 76638 7922 76690
rect 8878 76638 8930 76690
rect 9886 76638 9938 76690
rect 11006 76638 11058 76690
rect 43374 76638 43426 76690
rect 46734 76638 46786 76690
rect 47070 76638 47122 76690
rect 51662 76638 51714 76690
rect 55806 76638 55858 76690
rect 61294 76638 61346 76690
rect 61854 76638 61906 76690
rect 62526 76638 62578 76690
rect 63198 76638 63250 76690
rect 72382 76638 72434 76690
rect 73054 76638 73106 76690
rect 73950 76638 74002 76690
rect 74622 76638 74674 76690
rect 75294 76638 75346 76690
rect 76302 76638 76354 76690
rect 76974 76638 77026 76690
rect 77758 76638 77810 76690
rect 1934 76526 1986 76578
rect 5854 76526 5906 76578
rect 11678 76526 11730 76578
rect 13806 76526 13858 76578
rect 17726 76526 17778 76578
rect 29486 76526 29538 76578
rect 30158 76526 30210 76578
rect 32398 76526 32450 76578
rect 37214 76526 37266 76578
rect 38110 76526 38162 76578
rect 38894 76526 38946 76578
rect 42030 76526 42082 76578
rect 44942 76526 44994 76578
rect 45278 76526 45330 76578
rect 45838 76526 45890 76578
rect 47742 76526 47794 76578
rect 48078 76526 48130 76578
rect 48974 76526 49026 76578
rect 49870 76526 49922 76578
rect 50094 76526 50146 76578
rect 50766 76526 50818 76578
rect 50990 76526 51042 76578
rect 54798 76526 54850 76578
rect 57934 76526 57986 76578
rect 58942 76526 58994 76578
rect 59278 76526 59330 76578
rect 60958 76526 61010 76578
rect 64430 76526 64482 76578
rect 67230 76526 67282 76578
rect 70590 76526 70642 76578
rect 71486 76526 71538 76578
rect 6862 76414 6914 76466
rect 12798 76414 12850 76466
rect 14926 76414 14978 76466
rect 16718 76414 16770 76466
rect 18846 76414 18898 76466
rect 20638 76414 20690 76466
rect 22766 76414 22818 76466
rect 24558 76414 24610 76466
rect 26574 76414 26626 76466
rect 28478 76414 28530 76466
rect 31054 76414 31106 76466
rect 32174 76414 32226 76466
rect 33294 76414 33346 76466
rect 35086 76414 35138 76466
rect 37102 76414 37154 76466
rect 43038 76414 43090 76466
rect 43262 76414 43314 76466
rect 43486 76414 43538 76466
rect 43598 76414 43650 76466
rect 46174 76414 46226 76466
rect 49086 76414 49138 76466
rect 49646 76414 49698 76466
rect 51102 76414 51154 76466
rect 51998 76414 52050 76466
rect 63758 76414 63810 76466
rect 73278 76414 73330 76466
rect 3278 76302 3330 76354
rect 15710 76302 15762 76354
rect 19630 76302 19682 76354
rect 21870 76302 21922 76354
rect 23774 76302 23826 76354
rect 25790 76302 25842 76354
rect 27806 76302 27858 76354
rect 33966 76302 34018 76354
rect 35870 76302 35922 76354
rect 37886 76302 37938 76354
rect 40238 76302 40290 76354
rect 41022 76302 41074 76354
rect 44270 76302 44322 76354
rect 49982 76302 50034 76354
rect 56926 76302 56978 76354
rect 59726 76302 59778 76354
rect 37214 76190 37266 76242
rect 38222 76190 38274 76242
rect 48974 76190 49026 76242
rect 52670 76190 52722 76242
rect 64878 76190 64930 76242
rect 68350 76190 68402 76242
rect 4478 76022 4530 76074
rect 4582 76022 4634 76074
rect 4686 76022 4738 76074
rect 35198 76022 35250 76074
rect 35302 76022 35354 76074
rect 35406 76022 35458 76074
rect 65918 76022 65970 76074
rect 66022 76022 66074 76074
rect 66126 76022 66178 76074
rect 1822 75742 1874 75794
rect 7870 75742 7922 75794
rect 19854 75742 19906 75794
rect 20862 75742 20914 75794
rect 23998 75742 24050 75794
rect 24782 75742 24834 75794
rect 32734 75742 32786 75794
rect 36206 75742 36258 75794
rect 12910 75630 12962 75682
rect 15822 75630 15874 75682
rect 17838 75630 17890 75682
rect 26574 75630 26626 75682
rect 30158 75630 30210 75682
rect 30382 75630 30434 75682
rect 30942 75630 30994 75682
rect 31278 75630 31330 75682
rect 31502 75630 31554 75682
rect 32062 75630 32114 75682
rect 36094 75630 36146 75682
rect 5854 75518 5906 75570
rect 7198 75518 7250 75570
rect 13694 75518 13746 75570
rect 15262 75518 15314 75570
rect 17278 75518 17330 75570
rect 19294 75518 19346 75570
rect 21646 75518 21698 75570
rect 23326 75518 23378 75570
rect 25342 75518 25394 75570
rect 27134 75518 27186 75570
rect 27918 75518 27970 75570
rect 28478 75518 28530 75570
rect 28814 75518 28866 75570
rect 29822 75518 29874 75570
rect 33854 75518 33906 75570
rect 34078 75518 34130 75570
rect 34302 75518 34354 75570
rect 34414 75518 34466 75570
rect 35198 75518 35250 75570
rect 35534 75518 35586 75570
rect 36766 75518 36818 75570
rect 36318 75406 36370 75458
rect 37886 75854 37938 75906
rect 40910 75854 40962 75906
rect 41582 75854 41634 75906
rect 43486 75854 43538 75906
rect 46734 75854 46786 75906
rect 57262 75854 57314 75906
rect 70926 75854 70978 75906
rect 38782 75742 38834 75794
rect 40462 75742 40514 75794
rect 46286 75742 46338 75794
rect 49758 75742 49810 75794
rect 50878 75742 50930 75794
rect 52558 75742 52610 75794
rect 54126 75742 54178 75794
rect 56366 75742 56418 75794
rect 56926 75742 56978 75794
rect 62862 75742 62914 75794
rect 68686 75742 68738 75794
rect 38110 75630 38162 75682
rect 40686 75630 40738 75682
rect 43038 75630 43090 75682
rect 50766 75630 50818 75682
rect 50990 75630 51042 75682
rect 51774 75630 51826 75682
rect 52222 75630 52274 75682
rect 54350 75630 54402 75682
rect 61294 75630 61346 75682
rect 61630 75630 61682 75682
rect 62190 75630 62242 75682
rect 73950 75630 74002 75682
rect 40014 75518 40066 75570
rect 41806 75518 41858 75570
rect 42814 75518 42866 75570
rect 42926 75518 42978 75570
rect 44382 75518 44434 75570
rect 45838 75518 45890 75570
rect 48862 75518 48914 75570
rect 53678 75518 53730 75570
rect 55022 75518 55074 75570
rect 58158 75518 58210 75570
rect 59950 75518 60002 75570
rect 60510 75518 60562 75570
rect 62302 75518 62354 75570
rect 64990 75518 65042 75570
rect 66670 75518 66722 75570
rect 68014 75518 68066 75570
rect 69358 75518 69410 75570
rect 70254 75518 70306 75570
rect 73054 75518 73106 75570
rect 76078 75518 76130 75570
rect 77198 75518 77250 75570
rect 78094 75518 78146 75570
rect 36542 75406 36594 75458
rect 37326 75406 37378 75458
rect 37662 75406 37714 75458
rect 40126 75406 40178 75458
rect 40238 75406 40290 75458
rect 41246 75406 41298 75458
rect 42142 75406 42194 75458
rect 44046 75406 44098 75458
rect 45502 75406 45554 75458
rect 50542 75406 50594 75458
rect 51550 75406 51602 75458
rect 51662 75406 51714 75458
rect 53790 75406 53842 75458
rect 53902 75406 53954 75458
rect 57038 75406 57090 75458
rect 57822 75406 57874 75458
rect 58718 75406 58770 75458
rect 59054 75406 59106 75458
rect 59614 75406 59666 75458
rect 61518 75406 61570 75458
rect 65998 75406 66050 75458
rect 67342 75406 67394 75458
rect 69694 75406 69746 75458
rect 19838 75238 19890 75290
rect 19942 75238 19994 75290
rect 20046 75238 20098 75290
rect 50558 75238 50610 75290
rect 50662 75238 50714 75290
rect 50766 75238 50818 75290
rect 28142 75070 28194 75122
rect 29038 75070 29090 75122
rect 30270 75070 30322 75122
rect 30942 75070 30994 75122
rect 32286 75070 32338 75122
rect 34302 75070 34354 75122
rect 35310 75070 35362 75122
rect 36542 75070 36594 75122
rect 39454 75070 39506 75122
rect 39678 75070 39730 75122
rect 39790 75070 39842 75122
rect 40798 75070 40850 75122
rect 41694 75070 41746 75122
rect 41806 75070 41858 75122
rect 44270 75070 44322 75122
rect 44718 75070 44770 75122
rect 46734 75070 46786 75122
rect 47518 75070 47570 75122
rect 50094 75070 50146 75122
rect 54238 75070 54290 75122
rect 55358 75070 55410 75122
rect 57598 75070 57650 75122
rect 60622 75070 60674 75122
rect 61966 75070 62018 75122
rect 62638 75070 62690 75122
rect 63310 75070 63362 75122
rect 63982 75070 64034 75122
rect 65438 75070 65490 75122
rect 68350 75070 68402 75122
rect 69134 75070 69186 75122
rect 70814 75070 70866 75122
rect 73278 75070 73330 75122
rect 31166 74958 31218 75010
rect 33742 74958 33794 75010
rect 37438 74958 37490 75010
rect 38782 74958 38834 75010
rect 40462 74958 40514 75010
rect 45502 74958 45554 75010
rect 46846 74958 46898 75010
rect 48638 74958 48690 75010
rect 49982 74958 50034 75010
rect 50318 74958 50370 75010
rect 53006 74958 53058 75010
rect 54126 74958 54178 75010
rect 55246 74958 55298 75010
rect 56366 74958 56418 75010
rect 56702 74958 56754 75010
rect 58158 74958 58210 75010
rect 58718 74958 58770 75010
rect 60734 74958 60786 75010
rect 77646 74958 77698 75010
rect 29374 74846 29426 74898
rect 30046 74846 30098 74898
rect 30718 74846 30770 74898
rect 31278 74846 31330 74898
rect 32846 74846 32898 74898
rect 34190 74846 34242 74898
rect 34526 74846 34578 74898
rect 34638 74846 34690 74898
rect 37662 74846 37714 74898
rect 38446 74846 38498 74898
rect 39902 74846 39954 74898
rect 41582 74846 41634 74898
rect 42702 74846 42754 74898
rect 42926 74846 42978 74898
rect 43486 74846 43538 74898
rect 44158 74846 44210 74898
rect 44494 74846 44546 74898
rect 44718 74846 44770 74898
rect 45726 74846 45778 74898
rect 46174 74846 46226 74898
rect 46510 74846 46562 74898
rect 47854 74846 47906 74898
rect 48526 74846 48578 74898
rect 49534 74846 49586 74898
rect 51662 74846 51714 74898
rect 53230 74846 53282 74898
rect 53902 74846 53954 74898
rect 54350 74846 54402 74898
rect 54686 74846 54738 74898
rect 55470 74846 55522 74898
rect 55918 74846 55970 74898
rect 59390 74846 59442 74898
rect 59614 74846 59666 74898
rect 59950 74846 60002 74898
rect 61406 74846 61458 74898
rect 28590 74734 28642 74786
rect 32622 74734 32674 74786
rect 35870 74734 35922 74786
rect 42814 74734 42866 74786
rect 45614 74734 45666 74786
rect 49982 74734 50034 74786
rect 51214 74734 51266 74786
rect 52110 74734 52162 74786
rect 59502 74734 59554 74786
rect 64542 74734 64594 74786
rect 35646 74622 35698 74674
rect 36878 74622 36930 74674
rect 43262 74622 43314 74674
rect 57934 74622 57986 74674
rect 60622 74622 60674 74674
rect 61294 74622 61346 74674
rect 74510 74622 74562 74674
rect 4478 74454 4530 74506
rect 4582 74454 4634 74506
rect 4686 74454 4738 74506
rect 35198 74454 35250 74506
rect 35302 74454 35354 74506
rect 35406 74454 35458 74506
rect 65918 74454 65970 74506
rect 66022 74454 66074 74506
rect 66126 74454 66178 74506
rect 32286 74286 32338 74338
rect 33070 74286 33122 74338
rect 34190 74286 34242 74338
rect 44270 74286 44322 74338
rect 44382 74286 44434 74338
rect 45726 74286 45778 74338
rect 48414 74286 48466 74338
rect 49758 74286 49810 74338
rect 51662 74286 51714 74338
rect 56142 74286 56194 74338
rect 57038 74286 57090 74338
rect 59838 74286 59890 74338
rect 28814 74174 28866 74226
rect 29710 74174 29762 74226
rect 32174 74174 32226 74226
rect 32846 74174 32898 74226
rect 34526 74174 34578 74226
rect 37998 74174 38050 74226
rect 40126 74174 40178 74226
rect 42142 74174 42194 74226
rect 42702 74174 42754 74226
rect 44046 74174 44098 74226
rect 45950 74174 46002 74226
rect 48526 74174 48578 74226
rect 54014 74174 54066 74226
rect 54238 74174 54290 74226
rect 56366 74174 56418 74226
rect 57374 74174 57426 74226
rect 61966 74174 62018 74226
rect 62414 74174 62466 74226
rect 62862 74174 62914 74226
rect 63310 74174 63362 74226
rect 78094 74174 78146 74226
rect 31950 74062 32002 74114
rect 34750 74062 34802 74114
rect 35310 74062 35362 74114
rect 35534 74062 35586 74114
rect 35982 74062 36034 74114
rect 36542 74062 36594 74114
rect 36878 74062 36930 74114
rect 37550 74062 37602 74114
rect 38894 74062 38946 74114
rect 39566 74062 39618 74114
rect 40574 74062 40626 74114
rect 40686 74062 40738 74114
rect 40798 74062 40850 74114
rect 41246 74062 41298 74114
rect 42030 74062 42082 74114
rect 43038 74062 43090 74114
rect 43934 74062 43986 74114
rect 46174 74062 46226 74114
rect 46398 74062 46450 74114
rect 50542 74062 50594 74114
rect 51102 74062 51154 74114
rect 52222 74062 52274 74114
rect 52558 74062 52610 74114
rect 53454 74062 53506 74114
rect 54462 74062 54514 74114
rect 55470 74062 55522 74114
rect 55918 74062 55970 74114
rect 59166 74062 59218 74114
rect 59390 74062 59442 74114
rect 59614 74062 59666 74114
rect 60286 74062 60338 74114
rect 30158 73950 30210 74002
rect 30494 73950 30546 74002
rect 31054 73950 31106 74002
rect 35422 73950 35474 74002
rect 37998 73950 38050 74002
rect 38110 73950 38162 74002
rect 39006 73950 39058 74002
rect 42254 73950 42306 74002
rect 50206 73950 50258 74002
rect 50318 73950 50370 74002
rect 51326 73950 51378 74002
rect 51774 73950 51826 74002
rect 53566 73950 53618 74002
rect 57262 73950 57314 74002
rect 57934 73950 57986 74002
rect 58270 73950 58322 74002
rect 60622 73950 60674 74002
rect 31390 73838 31442 73890
rect 33406 73838 33458 73890
rect 36654 73838 36706 73890
rect 38334 73838 38386 73890
rect 39118 73838 39170 73890
rect 46286 73838 46338 73890
rect 47070 73838 47122 73890
rect 47742 73838 47794 73890
rect 49086 73838 49138 73890
rect 51550 73838 51602 73890
rect 52446 73838 52498 73890
rect 58046 73838 58098 73890
rect 59278 73838 59330 73890
rect 60510 73838 60562 73890
rect 61406 73838 61458 73890
rect 19838 73670 19890 73722
rect 19942 73670 19994 73722
rect 20046 73670 20098 73722
rect 50558 73670 50610 73722
rect 50662 73670 50714 73722
rect 50766 73670 50818 73722
rect 29486 73502 29538 73554
rect 30494 73502 30546 73554
rect 31390 73502 31442 73554
rect 32062 73502 32114 73554
rect 32958 73502 33010 73554
rect 33630 73502 33682 73554
rect 34862 73502 34914 73554
rect 35758 73502 35810 73554
rect 36430 73502 36482 73554
rect 40238 73502 40290 73554
rect 40350 73502 40402 73554
rect 40574 73502 40626 73554
rect 41470 73502 41522 73554
rect 41694 73502 41746 73554
rect 43822 73502 43874 73554
rect 47518 73502 47570 73554
rect 50542 73502 50594 73554
rect 55470 73502 55522 73554
rect 56142 73502 56194 73554
rect 56254 73502 56306 73554
rect 57598 73502 57650 73554
rect 60846 73502 60898 73554
rect 61406 73502 61458 73554
rect 61854 73502 61906 73554
rect 62302 73502 62354 73554
rect 62862 73502 62914 73554
rect 31278 73390 31330 73442
rect 31502 73390 31554 73442
rect 34526 73390 34578 73442
rect 37550 73390 37602 73442
rect 40798 73390 40850 73442
rect 41806 73390 41858 73442
rect 45390 73390 45442 73442
rect 48526 73390 48578 73442
rect 48750 73390 48802 73442
rect 51102 73390 51154 73442
rect 51774 73390 51826 73442
rect 52782 73390 52834 73442
rect 54462 73390 54514 73442
rect 57822 73390 57874 73442
rect 60286 73390 60338 73442
rect 33854 73278 33906 73330
rect 37438 73278 37490 73330
rect 38222 73278 38274 73330
rect 38670 73278 38722 73330
rect 44606 73278 44658 73330
rect 45278 73278 45330 73330
rect 46398 73278 46450 73330
rect 51886 73278 51938 73330
rect 52558 73278 52610 73330
rect 53566 73278 53618 73330
rect 54574 73278 54626 73330
rect 54798 73278 54850 73330
rect 56030 73278 56082 73330
rect 56702 73278 56754 73330
rect 59054 73278 59106 73330
rect 29934 73166 29986 73218
rect 30382 73166 30434 73218
rect 39118 73166 39170 73218
rect 39790 73166 39842 73218
rect 42590 73166 42642 73218
rect 45950 73166 46002 73218
rect 46286 73166 46338 73218
rect 48638 73166 48690 73218
rect 49646 73166 49698 73218
rect 52110 73166 52162 73218
rect 58606 73166 58658 73218
rect 59390 73166 59442 73218
rect 36766 73054 36818 73106
rect 42814 73054 42866 73106
rect 43038 73054 43090 73106
rect 43486 73054 43538 73106
rect 44830 73054 44882 73106
rect 45278 73054 45330 73106
rect 49870 73054 49922 73106
rect 50094 73054 50146 73106
rect 50990 73054 51042 73106
rect 54910 73054 54962 73106
rect 57486 73054 57538 73106
rect 60174 73054 60226 73106
rect 4478 72886 4530 72938
rect 4582 72886 4634 72938
rect 4686 72886 4738 72938
rect 35198 72886 35250 72938
rect 35302 72886 35354 72938
rect 35406 72886 35458 72938
rect 65918 72886 65970 72938
rect 66022 72886 66074 72938
rect 66126 72886 66178 72938
rect 36654 72718 36706 72770
rect 47070 72718 47122 72770
rect 57150 72718 57202 72770
rect 59614 72718 59666 72770
rect 60174 72718 60226 72770
rect 30942 72606 30994 72658
rect 32622 72606 32674 72658
rect 33070 72606 33122 72658
rect 33406 72606 33458 72658
rect 33854 72606 33906 72658
rect 43150 72606 43202 72658
rect 43934 72606 43986 72658
rect 47182 72606 47234 72658
rect 52446 72606 52498 72658
rect 54350 72606 54402 72658
rect 55806 72606 55858 72658
rect 56590 72606 56642 72658
rect 59390 72606 59442 72658
rect 59838 72606 59890 72658
rect 60286 72606 60338 72658
rect 61294 72606 61346 72658
rect 35086 72494 35138 72546
rect 37774 72494 37826 72546
rect 39118 72494 39170 72546
rect 40126 72494 40178 72546
rect 41582 72494 41634 72546
rect 42702 72494 42754 72546
rect 44046 72494 44098 72546
rect 44494 72494 44546 72546
rect 45614 72494 45666 72546
rect 46174 72494 46226 72546
rect 49870 72494 49922 72546
rect 50094 72494 50146 72546
rect 50430 72494 50482 72546
rect 52110 72494 52162 72546
rect 52670 72494 52722 72546
rect 53454 72494 53506 72546
rect 53902 72494 53954 72546
rect 55358 72494 55410 72546
rect 57038 72494 57090 72546
rect 57486 72494 57538 72546
rect 57822 72494 57874 72546
rect 58046 72494 58098 72546
rect 59278 72494 59330 72546
rect 34414 72382 34466 72434
rect 34526 72382 34578 72434
rect 35198 72382 35250 72434
rect 35982 72382 36034 72434
rect 36542 72382 36594 72434
rect 36654 72382 36706 72434
rect 37438 72382 37490 72434
rect 38894 72382 38946 72434
rect 41694 72382 41746 72434
rect 42254 72382 42306 72434
rect 45502 72382 45554 72434
rect 47742 72382 47794 72434
rect 48414 72382 48466 72434
rect 49310 72382 49362 72434
rect 55022 72382 55074 72434
rect 31950 72270 32002 72322
rect 37662 72270 37714 72322
rect 40238 72270 40290 72322
rect 41470 72270 41522 72322
rect 43822 72270 43874 72322
rect 49982 72270 50034 72322
rect 50878 72270 50930 72322
rect 19838 72102 19890 72154
rect 19942 72102 19994 72154
rect 20046 72102 20098 72154
rect 50558 72102 50610 72154
rect 50662 72102 50714 72154
rect 50766 72102 50818 72154
rect 33966 71934 34018 71986
rect 34302 71934 34354 71986
rect 35422 71934 35474 71986
rect 36094 71934 36146 71986
rect 36430 71934 36482 71986
rect 37102 71934 37154 71986
rect 37998 71934 38050 71986
rect 41470 71934 41522 71986
rect 43598 71934 43650 71986
rect 44942 71934 44994 71986
rect 45166 71934 45218 71986
rect 45950 71934 46002 71986
rect 46622 71934 46674 71986
rect 47294 71934 47346 71986
rect 47742 71934 47794 71986
rect 48638 71934 48690 71986
rect 53902 71934 53954 71986
rect 56590 71934 56642 71986
rect 59054 71934 59106 71986
rect 59614 71934 59666 71986
rect 34750 71822 34802 71874
rect 36990 71822 37042 71874
rect 43486 71822 43538 71874
rect 44158 71822 44210 71874
rect 46062 71822 46114 71874
rect 49758 71822 49810 71874
rect 52446 71822 52498 71874
rect 52782 71822 52834 71874
rect 55470 71822 55522 71874
rect 58606 71822 58658 71874
rect 37774 71710 37826 71762
rect 38782 71710 38834 71762
rect 39118 71710 39170 71762
rect 40462 71710 40514 71762
rect 42142 71710 42194 71762
rect 43038 71710 43090 71762
rect 43822 71710 43874 71762
rect 45278 71710 45330 71762
rect 45726 71710 45778 71762
rect 50318 71710 50370 71762
rect 51326 71710 51378 71762
rect 52558 71710 52610 71762
rect 52894 71710 52946 71762
rect 54238 71710 54290 71762
rect 54462 71710 54514 71762
rect 55246 71710 55298 71762
rect 56030 71710 56082 71762
rect 58046 71710 58098 71762
rect 39230 71598 39282 71650
rect 40350 71598 40402 71650
rect 48190 71598 48242 71650
rect 51774 71598 51826 71650
rect 57822 71598 57874 71650
rect 40238 71486 40290 71538
rect 48190 71486 48242 71538
rect 48638 71486 48690 71538
rect 56254 71486 56306 71538
rect 4478 71318 4530 71370
rect 4582 71318 4634 71370
rect 4686 71318 4738 71370
rect 35198 71318 35250 71370
rect 35302 71318 35354 71370
rect 35406 71318 35458 71370
rect 65918 71318 65970 71370
rect 66022 71318 66074 71370
rect 66126 71318 66178 71370
rect 33630 71150 33682 71202
rect 34750 71150 34802 71202
rect 39118 71150 39170 71202
rect 39678 71150 39730 71202
rect 40014 71150 40066 71202
rect 49198 71150 49250 71202
rect 50318 71150 50370 71202
rect 54462 71150 54514 71202
rect 54686 71150 54738 71202
rect 55022 71150 55074 71202
rect 55246 71150 55298 71202
rect 34750 71038 34802 71090
rect 35310 71038 35362 71090
rect 36430 71038 36482 71090
rect 36878 71038 36930 71090
rect 37662 71038 37714 71090
rect 38558 71038 38610 71090
rect 41022 71038 41074 71090
rect 42366 71038 42418 71090
rect 44158 71038 44210 71090
rect 45390 71038 45442 71090
rect 45950 71038 46002 71090
rect 46734 71038 46786 71090
rect 47406 71038 47458 71090
rect 47854 71038 47906 71090
rect 48302 71038 48354 71090
rect 49198 71038 49250 71090
rect 49758 71038 49810 71090
rect 50318 71038 50370 71090
rect 50878 71038 50930 71090
rect 54686 71038 54738 71090
rect 55246 71038 55298 71090
rect 55694 71038 55746 71090
rect 58942 71038 58994 71090
rect 38782 70926 38834 70978
rect 39678 70926 39730 70978
rect 41246 70926 41298 70978
rect 41806 70926 41858 70978
rect 42814 70926 42866 70978
rect 44494 70926 44546 70978
rect 48750 70926 48802 70978
rect 57038 70926 57090 70978
rect 38110 70814 38162 70866
rect 51550 70814 51602 70866
rect 52222 70814 52274 70866
rect 53566 70814 53618 70866
rect 56926 70814 56978 70866
rect 58270 70814 58322 70866
rect 46286 70702 46338 70754
rect 54126 70702 54178 70754
rect 58158 70702 58210 70754
rect 19838 70534 19890 70586
rect 19942 70534 19994 70586
rect 20046 70534 20098 70586
rect 50558 70534 50610 70586
rect 50662 70534 50714 70586
rect 50766 70534 50818 70586
rect 37102 70366 37154 70418
rect 37998 70366 38050 70418
rect 39006 70366 39058 70418
rect 39566 70366 39618 70418
rect 41582 70366 41634 70418
rect 42702 70366 42754 70418
rect 43598 70366 43650 70418
rect 44718 70366 44770 70418
rect 45054 70366 45106 70418
rect 45502 70366 45554 70418
rect 46398 70366 46450 70418
rect 46846 70366 46898 70418
rect 47182 70366 47234 70418
rect 48414 70366 48466 70418
rect 50430 70366 50482 70418
rect 51326 70366 51378 70418
rect 51774 70366 51826 70418
rect 52222 70366 52274 70418
rect 52670 70366 52722 70418
rect 53118 70366 53170 70418
rect 53566 70366 53618 70418
rect 54574 70366 54626 70418
rect 55022 70366 55074 70418
rect 55582 70366 55634 70418
rect 56366 70366 56418 70418
rect 37438 70254 37490 70306
rect 39678 70254 39730 70306
rect 40350 70254 40402 70306
rect 40798 70254 40850 70306
rect 43038 70254 43090 70306
rect 55470 70254 55522 70306
rect 40238 70142 40290 70194
rect 42366 70142 42418 70194
rect 42814 70142 42866 70194
rect 43934 70142 43986 70194
rect 44158 70142 44210 70194
rect 38334 70030 38386 70082
rect 37550 69918 37602 69970
rect 38334 69918 38386 69970
rect 4478 69750 4530 69802
rect 4582 69750 4634 69802
rect 4686 69750 4738 69802
rect 35198 69750 35250 69802
rect 35302 69750 35354 69802
rect 35406 69750 35458 69802
rect 65918 69750 65970 69802
rect 66022 69750 66074 69802
rect 66126 69750 66178 69802
rect 38334 69582 38386 69634
rect 39790 69582 39842 69634
rect 39790 69470 39842 69522
rect 40350 69470 40402 69522
rect 40798 69470 40850 69522
rect 46174 69470 46226 69522
rect 46622 69470 46674 69522
rect 52334 69470 52386 69522
rect 52782 69470 52834 69522
rect 19838 68966 19890 69018
rect 19942 68966 19994 69018
rect 20046 68966 20098 69018
rect 50558 68966 50610 69018
rect 50662 68966 50714 69018
rect 50766 68966 50818 69018
rect 4478 68182 4530 68234
rect 4582 68182 4634 68234
rect 4686 68182 4738 68234
rect 35198 68182 35250 68234
rect 35302 68182 35354 68234
rect 35406 68182 35458 68234
rect 65918 68182 65970 68234
rect 66022 68182 66074 68234
rect 66126 68182 66178 68234
rect 19838 67398 19890 67450
rect 19942 67398 19994 67450
rect 20046 67398 20098 67450
rect 50558 67398 50610 67450
rect 50662 67398 50714 67450
rect 50766 67398 50818 67450
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 35198 66614 35250 66666
rect 35302 66614 35354 66666
rect 35406 66614 35458 66666
rect 65918 66614 65970 66666
rect 66022 66614 66074 66666
rect 66126 66614 66178 66666
rect 19838 65830 19890 65882
rect 19942 65830 19994 65882
rect 20046 65830 20098 65882
rect 50558 65830 50610 65882
rect 50662 65830 50714 65882
rect 50766 65830 50818 65882
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 35198 65046 35250 65098
rect 35302 65046 35354 65098
rect 35406 65046 35458 65098
rect 65918 65046 65970 65098
rect 66022 65046 66074 65098
rect 66126 65046 66178 65098
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 50558 64262 50610 64314
rect 50662 64262 50714 64314
rect 50766 64262 50818 64314
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 65918 63478 65970 63530
rect 66022 63478 66074 63530
rect 66126 63478 66178 63530
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 50558 62694 50610 62746
rect 50662 62694 50714 62746
rect 50766 62694 50818 62746
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 65918 61910 65970 61962
rect 66022 61910 66074 61962
rect 66126 61910 66178 61962
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 50558 61126 50610 61178
rect 50662 61126 50714 61178
rect 50766 61126 50818 61178
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 65918 60342 65970 60394
rect 66022 60342 66074 60394
rect 66126 60342 66178 60394
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 50558 59558 50610 59610
rect 50662 59558 50714 59610
rect 50766 59558 50818 59610
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 65918 58774 65970 58826
rect 66022 58774 66074 58826
rect 66126 58774 66178 58826
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 50558 57990 50610 58042
rect 50662 57990 50714 58042
rect 50766 57990 50818 58042
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 65918 57206 65970 57258
rect 66022 57206 66074 57258
rect 66126 57206 66178 57258
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 65918 55638 65970 55690
rect 66022 55638 66074 55690
rect 66126 55638 66178 55690
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 65918 54070 65970 54122
rect 66022 54070 66074 54122
rect 66126 54070 66178 54122
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 65918 52502 65970 52554
rect 66022 52502 66074 52554
rect 66126 52502 66178 52554
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 65918 50934 65970 50986
rect 66022 50934 66074 50986
rect 66126 50934 66178 50986
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 65918 49366 65970 49418
rect 66022 49366 66074 49418
rect 66126 49366 66178 49418
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 65918 47798 65970 47850
rect 66022 47798 66074 47850
rect 66126 47798 66178 47850
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 65918 46230 65970 46282
rect 66022 46230 66074 46282
rect 66126 46230 66178 46282
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 65918 44662 65970 44714
rect 66022 44662 66074 44714
rect 66126 44662 66178 44714
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 65918 43094 65970 43146
rect 66022 43094 66074 43146
rect 66126 43094 66178 43146
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 65918 41526 65970 41578
rect 66022 41526 66074 41578
rect 66126 41526 66178 41578
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 65918 39958 65970 40010
rect 66022 39958 66074 40010
rect 66126 39958 66178 40010
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 65918 38390 65970 38442
rect 66022 38390 66074 38442
rect 66126 38390 66178 38442
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 65918 36822 65970 36874
rect 66022 36822 66074 36874
rect 66126 36822 66178 36874
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 65918 35254 65970 35306
rect 66022 35254 66074 35306
rect 66126 35254 66178 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 65918 33686 65970 33738
rect 66022 33686 66074 33738
rect 66126 33686 66178 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 65918 32118 65970 32170
rect 66022 32118 66074 32170
rect 66126 32118 66178 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 65918 30550 65970 30602
rect 66022 30550 66074 30602
rect 66126 30550 66178 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 65918 28982 65970 29034
rect 66022 28982 66074 29034
rect 66126 28982 66178 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 65918 27414 65970 27466
rect 66022 27414 66074 27466
rect 66126 27414 66178 27466
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 65918 25846 65970 25898
rect 66022 25846 66074 25898
rect 66126 25846 66178 25898
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 65918 24278 65970 24330
rect 66022 24278 66074 24330
rect 66126 24278 66178 24330
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 65918 22710 65970 22762
rect 66022 22710 66074 22762
rect 66126 22710 66178 22762
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 65918 21142 65970 21194
rect 66022 21142 66074 21194
rect 66126 21142 66178 21194
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 65918 19574 65970 19626
rect 66022 19574 66074 19626
rect 66126 19574 66178 19626
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 65918 18006 65970 18058
rect 66022 18006 66074 18058
rect 66126 18006 66178 18058
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 65918 16438 65970 16490
rect 66022 16438 66074 16490
rect 66126 16438 66178 16490
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 65918 14870 65970 14922
rect 66022 14870 66074 14922
rect 66126 14870 66178 14922
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 65918 13302 65970 13354
rect 66022 13302 66074 13354
rect 66126 13302 66178 13354
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 65918 11734 65970 11786
rect 66022 11734 66074 11786
rect 66126 11734 66178 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 65918 10166 65970 10218
rect 66022 10166 66074 10218
rect 66126 10166 66178 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 65918 8598 65970 8650
rect 66022 8598 66074 8650
rect 66126 8598 66178 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 65918 7030 65970 7082
rect 66022 7030 66074 7082
rect 66126 7030 66178 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 65918 5462 65970 5514
rect 66022 5462 66074 5514
rect 66126 5462 66178 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 13918 4398 13970 4450
rect 17950 4398 18002 4450
rect 24670 4398 24722 4450
rect 29374 4398 29426 4450
rect 32510 4398 32562 4450
rect 37214 4398 37266 4450
rect 51326 4398 51378 4450
rect 55358 4398 55410 4450
rect 59390 4398 59442 4450
rect 63422 4398 63474 4450
rect 70814 4398 70866 4450
rect 73390 4398 73442 4450
rect 74062 4398 74114 4450
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 65918 3894 65970 3946
rect 66022 3894 66074 3946
rect 66126 3894 66178 3946
rect 6974 3278 7026 3330
rect 8094 3278 8146 3330
rect 8878 3278 8930 3330
rect 9998 3278 10050 3330
rect 10782 3278 10834 3330
rect 11454 3278 11506 3330
rect 12126 3278 12178 3330
rect 12798 3278 12850 3330
rect 14030 3278 14082 3330
rect 14702 3278 14754 3330
rect 15374 3278 15426 3330
rect 16046 3278 16098 3330
rect 16718 3278 16770 3330
rect 17950 3278 18002 3330
rect 18622 3278 18674 3330
rect 19294 3278 19346 3330
rect 19966 3278 20018 3330
rect 20638 3278 20690 3330
rect 21758 3278 21810 3330
rect 22430 3278 22482 3330
rect 23102 3278 23154 3330
rect 23774 3278 23826 3330
rect 24558 3278 24610 3330
rect 25790 3278 25842 3330
rect 26462 3278 26514 3330
rect 27134 3278 27186 3330
rect 27806 3278 27858 3330
rect 28478 3278 28530 3330
rect 29710 3278 29762 3330
rect 30270 3278 30322 3330
rect 30942 3278 30994 3330
rect 31614 3278 31666 3330
rect 32398 3278 32450 3330
rect 33630 3278 33682 3330
rect 34302 3278 34354 3330
rect 34974 3278 35026 3330
rect 35646 3278 35698 3330
rect 36318 3278 36370 3330
rect 37550 3278 37602 3330
rect 38222 3278 38274 3330
rect 38894 3278 38946 3330
rect 39566 3278 39618 3330
rect 40238 3278 40290 3330
rect 41246 3278 41298 3330
rect 41918 3278 41970 3330
rect 42590 3278 42642 3330
rect 43262 3278 43314 3330
rect 43934 3278 43986 3330
rect 44942 3278 44994 3330
rect 45614 3278 45666 3330
rect 46286 3278 46338 3330
rect 46958 3278 47010 3330
rect 47630 3278 47682 3330
rect 48862 3278 48914 3330
rect 49534 3278 49586 3330
rect 50206 3278 50258 3330
rect 50878 3278 50930 3330
rect 51550 3278 51602 3330
rect 52782 3278 52834 3330
rect 53454 3278 53506 3330
rect 54126 3278 54178 3330
rect 54798 3278 54850 3330
rect 55470 3278 55522 3330
rect 56702 3278 56754 3330
rect 57374 3278 57426 3330
rect 58046 3278 58098 3330
rect 58718 3278 58770 3330
rect 59390 3278 59442 3330
rect 60622 3278 60674 3330
rect 61294 3278 61346 3330
rect 61966 3278 62018 3330
rect 62638 3278 62690 3330
rect 63310 3278 63362 3330
rect 64542 3278 64594 3330
rect 65214 3278 65266 3330
rect 65886 3278 65938 3330
rect 66558 3278 66610 3330
rect 67230 3278 67282 3330
rect 68462 3278 68514 3330
rect 69134 3278 69186 3330
rect 69806 3278 69858 3330
rect 70478 3278 70530 3330
rect 71150 3278 71202 3330
rect 72382 3278 72434 3330
rect 73054 3278 73106 3330
rect 73726 3278 73778 3330
rect 74398 3278 74450 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
rect 46398 1822 46450 1874
rect 46958 1822 47010 1874
rect 57822 1822 57874 1874
rect 58718 1822 58770 1874
rect 61182 1822 61234 1874
rect 61966 1822 62018 1874
rect 64654 1822 64706 1874
rect 65214 1822 65266 1874
rect 65886 1822 65938 1874
rect 66558 1822 66610 1874
rect 24558 1710 24610 1762
rect 25118 1710 25170 1762
rect 32398 1710 32450 1762
rect 32958 1710 33010 1762
rect 44382 1710 44434 1762
rect 44942 1710 44994 1762
rect 45726 1710 45778 1762
rect 46286 1710 46338 1762
rect 47070 1710 47122 1762
rect 47630 1710 47682 1762
rect 49086 1710 49138 1762
rect 50206 1710 50258 1762
rect 50430 1710 50482 1762
rect 51550 1710 51602 1762
rect 52446 1710 52498 1762
rect 53454 1710 53506 1762
rect 53790 1710 53842 1762
rect 54798 1710 54850 1762
rect 55806 1710 55858 1762
rect 56702 1710 56754 1762
rect 57150 1710 57202 1762
rect 58046 1710 58098 1762
rect 60510 1710 60562 1762
rect 61294 1710 61346 1762
rect 62526 1710 62578 1762
rect 63310 1710 63362 1762
rect 63870 1710 63922 1762
rect 64542 1710 64594 1762
rect 67230 1710 67282 1762
rect 68462 1710 68514 1762
rect 69246 1710 69298 1762
rect 70478 1710 70530 1762
rect 72606 1710 72658 1762
rect 73726 1710 73778 1762
<< metal2 >>
rect 1568 79200 1680 80000
rect 2240 79200 2352 80000
rect 2912 79200 3024 80000
rect 3584 79200 3696 80000
rect 4256 79200 4368 80000
rect 4928 79200 5040 80000
rect 5600 79200 5712 80000
rect 6272 79200 6384 80000
rect 6944 79200 7056 80000
rect 7616 79200 7728 80000
rect 8288 79200 8400 80000
rect 8960 79200 9072 80000
rect 9632 79200 9744 80000
rect 10304 79200 10416 80000
rect 10976 79200 11088 80000
rect 11648 79200 11760 80000
rect 12320 79200 12432 80000
rect 12992 79200 13104 80000
rect 13664 79200 13776 80000
rect 14336 79200 14448 80000
rect 15008 79200 15120 80000
rect 15680 79200 15792 80000
rect 16352 79200 16464 80000
rect 17024 79200 17136 80000
rect 17696 79200 17808 80000
rect 18368 79200 18480 80000
rect 19040 79200 19152 80000
rect 19712 79200 19824 80000
rect 20384 79200 20496 80000
rect 21056 79200 21168 80000
rect 21728 79200 21840 80000
rect 22400 79200 22512 80000
rect 23072 79200 23184 80000
rect 23744 79200 23856 80000
rect 24416 79200 24528 80000
rect 25088 79200 25200 80000
rect 25760 79200 25872 80000
rect 26432 79200 26544 80000
rect 27104 79200 27216 80000
rect 27776 79200 27888 80000
rect 28448 79200 28560 80000
rect 29120 79200 29232 80000
rect 29792 79200 29904 80000
rect 30464 79200 30576 80000
rect 31136 79200 31248 80000
rect 31808 79200 31920 80000
rect 32480 79200 32592 80000
rect 33152 79200 33264 80000
rect 33824 79200 33936 80000
rect 34496 79200 34608 80000
rect 35168 79200 35280 80000
rect 35840 79200 35952 80000
rect 36512 79200 36624 80000
rect 37184 79200 37296 80000
rect 37856 79200 37968 80000
rect 38528 79200 38640 80000
rect 39200 79200 39312 80000
rect 39872 79200 39984 80000
rect 40544 79200 40656 80000
rect 41216 79200 41328 80000
rect 41888 79200 42000 80000
rect 42560 79200 42672 80000
rect 43232 79200 43344 80000
rect 43904 79200 44016 80000
rect 44576 79200 44688 80000
rect 45248 79200 45360 80000
rect 45920 79200 46032 80000
rect 46592 79200 46704 80000
rect 47264 79200 47376 80000
rect 47936 79200 48048 80000
rect 48608 79200 48720 80000
rect 49280 79200 49392 80000
rect 49952 79200 50064 80000
rect 50624 79200 50736 80000
rect 51296 79200 51408 80000
rect 51968 79200 52080 80000
rect 52640 79200 52752 80000
rect 53312 79200 53424 80000
rect 53984 79200 54096 80000
rect 54656 79200 54768 80000
rect 55328 79200 55440 80000
rect 56000 79200 56112 80000
rect 56672 79200 56784 80000
rect 57344 79200 57456 80000
rect 58016 79200 58128 80000
rect 58688 79200 58800 80000
rect 59360 79200 59472 80000
rect 60032 79200 60144 80000
rect 60704 79200 60816 80000
rect 61376 79200 61488 80000
rect 62048 79200 62160 80000
rect 62720 79200 62832 80000
rect 63392 79200 63504 80000
rect 64064 79200 64176 80000
rect 64736 79200 64848 80000
rect 65408 79200 65520 80000
rect 66080 79200 66192 80000
rect 66752 79200 66864 80000
rect 67424 79200 67536 80000
rect 68096 79200 68208 80000
rect 68768 79200 68880 80000
rect 69440 79200 69552 80000
rect 70112 79200 70224 80000
rect 70784 79200 70896 80000
rect 71456 79200 71568 80000
rect 72128 79200 72240 80000
rect 72800 79200 72912 80000
rect 73472 79200 73584 80000
rect 74144 79200 74256 80000
rect 74816 79200 74928 80000
rect 75488 79200 75600 80000
rect 76160 79200 76272 80000
rect 76832 79200 76944 80000
rect 77504 79200 77616 80000
rect 78176 79200 78288 80000
rect 1596 76580 1652 79200
rect 2940 76692 2996 79200
rect 2940 76626 2996 76636
rect 1932 76580 1988 76590
rect 1596 76578 1988 76580
rect 1596 76526 1934 76578
rect 1986 76526 1988 76578
rect 1596 76524 1988 76526
rect 1820 75794 1876 76524
rect 1932 76514 1988 76524
rect 3612 76580 3668 79200
rect 3836 76692 3892 76702
rect 3836 76598 3892 76636
rect 4956 76690 5012 79200
rect 4956 76638 4958 76690
rect 5010 76638 5012 76690
rect 4956 76626 5012 76638
rect 3612 76514 3668 76524
rect 3276 76356 3332 76366
rect 3276 76354 3444 76356
rect 3276 76302 3278 76354
rect 3330 76302 3444 76354
rect 3276 76300 3444 76302
rect 3276 76290 3332 76300
rect 3388 75908 3444 76300
rect 4476 76076 4740 76086
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4476 76010 4740 76020
rect 3388 75842 3444 75852
rect 1820 75742 1822 75794
rect 1874 75742 1876 75794
rect 1820 75730 1876 75742
rect 5628 75572 5684 79200
rect 6860 76692 6916 76702
rect 5852 76580 5908 76590
rect 5852 76486 5908 76524
rect 6860 76466 6916 76636
rect 6860 76414 6862 76466
rect 6914 76414 6916 76466
rect 6860 76402 6916 76414
rect 5852 75572 5908 75582
rect 5628 75570 5908 75572
rect 5628 75518 5854 75570
rect 5906 75518 5908 75570
rect 5628 75516 5908 75518
rect 6972 75572 7028 79200
rect 7644 76692 7700 79200
rect 7868 76692 7924 76702
rect 7644 76690 7924 76692
rect 7644 76638 7870 76690
rect 7922 76638 7924 76690
rect 7644 76636 7924 76638
rect 7868 76626 7924 76636
rect 7980 76692 8036 76702
rect 7868 75796 7924 75806
rect 7980 75796 8036 76636
rect 8876 76692 8932 76702
rect 8988 76692 9044 79200
rect 8876 76690 9044 76692
rect 8876 76638 8878 76690
rect 8930 76638 9044 76690
rect 8876 76636 9044 76638
rect 9660 76692 9716 79200
rect 9884 76692 9940 76702
rect 9660 76690 9940 76692
rect 9660 76638 9886 76690
rect 9938 76638 9940 76690
rect 9660 76636 9940 76638
rect 8876 76626 8932 76636
rect 9884 76626 9940 76636
rect 11004 76690 11060 79200
rect 11004 76638 11006 76690
rect 11058 76638 11060 76690
rect 11004 76626 11060 76638
rect 11676 76578 11732 79200
rect 11676 76526 11678 76578
rect 11730 76526 11732 76578
rect 11676 76514 11732 76526
rect 12796 76468 12852 76478
rect 12796 76466 12964 76468
rect 12796 76414 12798 76466
rect 12850 76414 12964 76466
rect 12796 76412 12964 76414
rect 12796 76402 12852 76412
rect 7868 75794 8036 75796
rect 7868 75742 7870 75794
rect 7922 75742 8036 75794
rect 7868 75740 8036 75742
rect 7868 75730 7924 75740
rect 12908 75682 12964 76412
rect 12908 75630 12910 75682
rect 12962 75630 12964 75682
rect 7196 75572 7252 75582
rect 6972 75570 7252 75572
rect 6972 75518 7198 75570
rect 7250 75518 7252 75570
rect 6972 75516 7252 75518
rect 5852 75506 5908 75516
rect 7196 75506 7252 75516
rect 4476 74508 4740 74518
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4476 74442 4740 74452
rect 4476 72940 4740 72950
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4476 72874 4740 72884
rect 12908 72548 12964 75630
rect 13020 75572 13076 79200
rect 13692 76580 13748 79200
rect 13804 76580 13860 76590
rect 13692 76578 13860 76580
rect 13692 76526 13806 76578
rect 13858 76526 13860 76578
rect 13692 76524 13860 76526
rect 13804 76514 13860 76524
rect 14924 76468 14980 76478
rect 14924 76374 14980 76412
rect 13020 75506 13076 75516
rect 13692 75572 13748 75582
rect 15036 75572 15092 79200
rect 15708 76354 15764 79200
rect 15708 76302 15710 76354
rect 15762 76302 15764 76354
rect 15708 76290 15764 76302
rect 15820 76468 15876 76478
rect 15820 75682 15876 76412
rect 15820 75630 15822 75682
rect 15874 75630 15876 75682
rect 15260 75572 15316 75582
rect 15036 75570 15316 75572
rect 15036 75518 15262 75570
rect 15314 75518 15316 75570
rect 15036 75516 15316 75518
rect 13692 75478 13748 75516
rect 15260 75506 15316 75516
rect 15820 75460 15876 75630
rect 16716 76466 16772 76478
rect 16716 76414 16718 76466
rect 16770 76414 16772 76466
rect 16716 75684 16772 76414
rect 16716 75618 16772 75628
rect 17052 75572 17108 79200
rect 17724 76578 17780 79200
rect 17724 76526 17726 76578
rect 17778 76526 17780 76578
rect 17724 76514 17780 76526
rect 18844 76468 18900 76478
rect 18844 76374 18900 76412
rect 17836 75684 17892 75694
rect 17836 75590 17892 75628
rect 17276 75572 17332 75582
rect 17052 75570 17332 75572
rect 17052 75518 17278 75570
rect 17330 75518 17332 75570
rect 17052 75516 17332 75518
rect 19068 75572 19124 79200
rect 19740 77812 19796 79200
rect 19628 77756 19796 77812
rect 19628 76354 19684 77756
rect 19836 76860 20100 76870
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 19836 76794 20100 76804
rect 19628 76302 19630 76354
rect 19682 76302 19684 76354
rect 19628 76290 19684 76302
rect 19852 76468 19908 76478
rect 19852 76244 19908 76412
rect 20636 76468 20692 76478
rect 20636 76466 20916 76468
rect 20636 76414 20638 76466
rect 20690 76414 20916 76466
rect 20636 76412 20916 76414
rect 20636 76402 20692 76412
rect 19852 75794 19908 76188
rect 19852 75742 19854 75794
rect 19906 75742 19908 75794
rect 19852 75730 19908 75742
rect 20860 76020 20916 76412
rect 20860 75794 20916 75964
rect 20860 75742 20862 75794
rect 20914 75742 20916 75794
rect 20860 75730 20916 75742
rect 19292 75572 19348 75582
rect 19068 75570 19348 75572
rect 19068 75518 19294 75570
rect 19346 75518 19348 75570
rect 19068 75516 19348 75518
rect 17276 75506 17332 75516
rect 19292 75506 19348 75516
rect 21084 75572 21140 79200
rect 21756 76356 21812 79200
rect 22764 76466 22820 76478
rect 22764 76414 22766 76466
rect 22818 76414 22820 76466
rect 21868 76356 21924 76366
rect 21756 76354 21924 76356
rect 21756 76302 21870 76354
rect 21922 76302 21924 76354
rect 21756 76300 21924 76302
rect 21868 76290 21924 76300
rect 21756 75908 21812 75918
rect 21084 75506 21140 75516
rect 21644 75572 21700 75582
rect 21644 75478 21700 75516
rect 15820 75394 15876 75404
rect 21420 75460 21476 75470
rect 19836 75292 20100 75302
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 19836 75226 20100 75236
rect 19836 73724 20100 73734
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 19836 73658 20100 73668
rect 12908 72482 12964 72492
rect 21420 72436 21476 75404
rect 21756 74340 21812 75852
rect 22764 75908 22820 76414
rect 22764 75842 22820 75852
rect 23100 75572 23156 79200
rect 23772 76354 23828 79200
rect 24556 76468 24612 76478
rect 24556 76466 24836 76468
rect 24556 76414 24558 76466
rect 24610 76414 24836 76466
rect 24556 76412 24836 76414
rect 24556 76402 24612 76412
rect 23772 76302 23774 76354
rect 23826 76302 23828 76354
rect 23772 76290 23828 76302
rect 23996 75908 24052 75918
rect 23996 75794 24052 75852
rect 23996 75742 23998 75794
rect 24050 75742 24052 75794
rect 23996 75730 24052 75742
rect 24780 75796 24836 76412
rect 24780 75664 24836 75740
rect 23324 75572 23380 75582
rect 23100 75570 23380 75572
rect 23100 75518 23326 75570
rect 23378 75518 23380 75570
rect 23100 75516 23380 75518
rect 25116 75572 25172 79200
rect 25788 76354 25844 79200
rect 25788 76302 25790 76354
rect 25842 76302 25844 76354
rect 25788 76290 25844 76302
rect 26572 76466 26628 76478
rect 26572 76414 26574 76466
rect 26626 76414 26628 76466
rect 26572 75682 26628 76414
rect 26572 75630 26574 75682
rect 26626 75630 26628 75682
rect 25340 75572 25396 75582
rect 25116 75570 25396 75572
rect 25116 75518 25342 75570
rect 25394 75518 25396 75570
rect 25116 75516 25396 75518
rect 23324 75506 23380 75516
rect 25340 75506 25396 75516
rect 26572 74452 26628 75630
rect 27132 75570 27188 79200
rect 27804 76354 27860 79200
rect 28476 76468 28532 76478
rect 28476 76466 28756 76468
rect 28476 76414 28478 76466
rect 28530 76414 28756 76466
rect 28476 76412 28756 76414
rect 28476 76402 28532 76412
rect 27804 76302 27806 76354
rect 27858 76302 27860 76354
rect 27804 76290 27860 76302
rect 28476 75796 28532 75806
rect 27132 75518 27134 75570
rect 27186 75518 27188 75570
rect 27132 75506 27188 75518
rect 27916 75572 27972 75582
rect 27916 75478 27972 75516
rect 28476 75570 28532 75740
rect 28476 75518 28478 75570
rect 28530 75518 28532 75570
rect 28140 75460 28196 75470
rect 28140 75122 28196 75404
rect 28140 75070 28142 75122
rect 28194 75070 28196 75122
rect 28140 75058 28196 75070
rect 26572 74386 26628 74396
rect 21756 74274 21812 74284
rect 28476 73444 28532 75518
rect 28700 75348 28756 76412
rect 29148 75796 29204 79200
rect 29820 77812 29876 79200
rect 29820 77756 30212 77812
rect 29484 76580 29540 76590
rect 29484 76578 29988 76580
rect 29484 76526 29486 76578
rect 29538 76526 29988 76578
rect 29484 76524 29988 76526
rect 29484 76514 29540 76524
rect 29148 75730 29204 75740
rect 28812 75572 28868 75582
rect 29820 75572 29876 75582
rect 28812 75570 29876 75572
rect 28812 75518 28814 75570
rect 28866 75518 29822 75570
rect 29874 75518 29876 75570
rect 28812 75516 29876 75518
rect 28812 75506 28868 75516
rect 29820 75506 29876 75516
rect 29932 75572 29988 76524
rect 30156 76578 30212 77756
rect 30156 76526 30158 76578
rect 30210 76526 30212 76578
rect 30156 76514 30212 76526
rect 31052 76468 31108 76478
rect 30604 76466 31108 76468
rect 30604 76414 31054 76466
rect 31106 76414 31108 76466
rect 30604 76412 31108 76414
rect 31164 76468 31220 79200
rect 31164 76412 31668 76468
rect 29932 75506 29988 75516
rect 30044 75684 30100 75694
rect 28700 75292 29092 75348
rect 29036 75122 29092 75292
rect 29036 75070 29038 75122
rect 29090 75070 29092 75122
rect 29036 75058 29092 75070
rect 29372 74898 29428 74910
rect 29372 74846 29374 74898
rect 29426 74846 29428 74898
rect 28588 74786 28644 74798
rect 28588 74734 28590 74786
rect 28642 74734 28644 74786
rect 28588 74228 28644 74734
rect 28588 74162 28644 74172
rect 28812 74340 28868 74350
rect 28812 74226 28868 74284
rect 29372 74340 29428 74846
rect 30044 74898 30100 75628
rect 30156 75682 30212 75694
rect 30156 75630 30158 75682
rect 30210 75630 30212 75682
rect 30156 75460 30212 75630
rect 30380 75684 30436 75694
rect 30380 75682 30548 75684
rect 30380 75630 30382 75682
rect 30434 75630 30548 75682
rect 30380 75628 30548 75630
rect 30380 75618 30436 75628
rect 30156 75394 30212 75404
rect 30492 75460 30548 75628
rect 30268 75124 30324 75134
rect 30268 75030 30324 75068
rect 30044 74846 30046 74898
rect 30098 74846 30100 74898
rect 30044 74834 30100 74846
rect 29372 74274 29428 74284
rect 28812 74174 28814 74226
rect 28866 74174 28868 74226
rect 28812 74004 28868 74174
rect 29708 74228 29764 74238
rect 29708 74134 29764 74172
rect 28812 73938 28868 73948
rect 29484 74004 29540 74014
rect 29484 73554 29540 73948
rect 30156 74004 30212 74014
rect 30156 73910 30212 73948
rect 30492 74002 30548 75404
rect 30492 73950 30494 74002
rect 30546 73950 30548 74002
rect 30492 73938 30548 73950
rect 29484 73502 29486 73554
rect 29538 73502 29540 73554
rect 29484 73490 29540 73502
rect 30492 73556 30548 73566
rect 30604 73556 30660 76412
rect 31052 76402 31108 76412
rect 30940 75684 30996 75694
rect 31276 75684 31332 75694
rect 30940 75590 30996 75628
rect 31164 75682 31332 75684
rect 31164 75630 31278 75682
rect 31330 75630 31332 75682
rect 31164 75628 31332 75630
rect 30716 75348 30772 75358
rect 30716 74900 30772 75292
rect 30940 75236 30996 75246
rect 30940 75122 30996 75180
rect 30940 75070 30942 75122
rect 30994 75070 30996 75122
rect 30940 75058 30996 75070
rect 31164 75236 31220 75628
rect 31276 75618 31332 75628
rect 31500 75682 31556 75694
rect 31500 75630 31502 75682
rect 31554 75630 31556 75682
rect 31500 75460 31556 75630
rect 31500 75394 31556 75404
rect 30716 74768 30772 74844
rect 31164 75010 31220 75180
rect 31164 74958 31166 75010
rect 31218 74958 31220 75010
rect 31164 74228 31220 74958
rect 31500 75124 31556 75134
rect 31164 74162 31220 74172
rect 31276 74898 31332 74910
rect 31276 74846 31278 74898
rect 31330 74846 31332 74898
rect 31052 74004 31108 74014
rect 31052 73910 31108 73948
rect 31276 73668 31332 74846
rect 31388 73892 31444 73902
rect 31388 73798 31444 73836
rect 31276 73612 31444 73668
rect 30492 73554 30660 73556
rect 30492 73502 30494 73554
rect 30546 73502 30660 73554
rect 30492 73500 30660 73502
rect 31388 73554 31444 73612
rect 31388 73502 31390 73554
rect 31442 73502 31444 73554
rect 30492 73490 30548 73500
rect 31388 73490 31444 73502
rect 28476 73378 28532 73388
rect 30940 73444 30996 73454
rect 29932 73220 29988 73230
rect 30380 73220 30436 73230
rect 29932 73218 30436 73220
rect 29932 73166 29934 73218
rect 29986 73166 30382 73218
rect 30434 73166 30436 73218
rect 29932 73164 30436 73166
rect 29932 73154 29988 73164
rect 30380 72772 30436 73164
rect 30380 72706 30436 72716
rect 30940 72658 30996 73388
rect 31276 73444 31332 73454
rect 31276 73350 31332 73388
rect 31500 73442 31556 75068
rect 31612 73556 31668 76412
rect 31836 75796 31892 79200
rect 32396 77026 32452 77038
rect 32396 76974 32398 77026
rect 32450 76974 32452 77026
rect 32396 76578 32452 76974
rect 32396 76526 32398 76578
rect 32450 76526 32452 76578
rect 31836 75730 31892 75740
rect 32172 76466 32228 76478
rect 32172 76414 32174 76466
rect 32226 76414 32228 76466
rect 32060 75682 32116 75694
rect 32060 75630 32062 75682
rect 32114 75630 32116 75682
rect 32060 75124 32116 75630
rect 32172 75124 32228 76414
rect 32284 75124 32340 75134
rect 32172 75122 32340 75124
rect 32172 75070 32286 75122
rect 32338 75070 32340 75122
rect 32172 75068 32340 75070
rect 32060 75058 32116 75068
rect 32284 75058 32340 75068
rect 32060 74900 32116 74910
rect 31948 74452 32004 74462
rect 31948 74114 32004 74396
rect 31948 74062 31950 74114
rect 32002 74062 32004 74114
rect 31948 74050 32004 74062
rect 32060 73892 32116 74844
rect 32284 74340 32340 74350
rect 32396 74340 32452 76526
rect 32732 75796 32788 75806
rect 32732 75702 32788 75740
rect 33180 75572 33236 79200
rect 33292 77026 33348 77038
rect 33292 76974 33294 77026
rect 33346 76974 33348 77026
rect 33292 76466 33348 76974
rect 33292 76414 33294 76466
rect 33346 76414 33348 76466
rect 33292 76402 33348 76414
rect 33852 76356 33908 79200
rect 34412 77700 34468 77710
rect 33964 76356 34020 76366
rect 33852 76354 34020 76356
rect 33852 76302 33966 76354
rect 34018 76302 34020 76354
rect 33852 76300 34020 76302
rect 33964 76290 34020 76300
rect 34300 76244 34356 76254
rect 34188 76020 34244 76030
rect 33180 75506 33236 75516
rect 33852 75570 33908 75582
rect 33852 75518 33854 75570
rect 33906 75518 33908 75570
rect 32844 75460 32900 75470
rect 32844 74898 32900 75404
rect 32844 74846 32846 74898
rect 32898 74846 32900 74898
rect 32620 74788 32676 74798
rect 32620 74694 32676 74732
rect 32284 74338 32452 74340
rect 32284 74286 32286 74338
rect 32338 74286 32452 74338
rect 32284 74284 32452 74286
rect 32620 74452 32676 74462
rect 32284 74274 32340 74284
rect 32172 74228 32228 74238
rect 32172 74134 32228 74172
rect 31612 73490 31668 73500
rect 31948 73836 32116 73892
rect 31500 73390 31502 73442
rect 31554 73390 31556 73442
rect 31500 73378 31556 73390
rect 30940 72606 30942 72658
rect 30994 72606 30996 72658
rect 30940 72594 30996 72606
rect 21420 72370 21476 72380
rect 31948 72322 32004 73836
rect 32060 73556 32116 73566
rect 32060 73462 32116 73500
rect 32620 73556 32676 74396
rect 32844 74226 32900 74846
rect 32844 74174 32846 74226
rect 32898 74174 32900 74226
rect 32844 74162 32900 74174
rect 33068 75124 33124 75134
rect 33068 74338 33124 75068
rect 33740 75012 33796 75022
rect 33740 74918 33796 74956
rect 33068 74286 33070 74338
rect 33122 74286 33124 74338
rect 32620 72658 32676 73500
rect 32956 73668 33012 73678
rect 32956 73554 33012 73612
rect 32956 73502 32958 73554
rect 33010 73502 33012 73554
rect 32956 73490 33012 73502
rect 32620 72606 32622 72658
rect 32674 72606 32676 72658
rect 32620 72594 32676 72606
rect 33068 72660 33124 74286
rect 33852 74228 33908 75518
rect 34076 75570 34132 75582
rect 34076 75518 34078 75570
rect 34130 75518 34132 75570
rect 34076 74788 34132 75518
rect 34188 75124 34244 75964
rect 34300 75570 34356 76188
rect 34300 75518 34302 75570
rect 34354 75518 34356 75570
rect 34300 75506 34356 75518
rect 34412 75570 34468 77644
rect 35196 76692 35252 79200
rect 34412 75518 34414 75570
rect 34466 75518 34468 75570
rect 34300 75124 34356 75134
rect 34188 75122 34356 75124
rect 34188 75070 34302 75122
rect 34354 75070 34356 75122
rect 34188 75068 34356 75070
rect 34300 75058 34356 75068
rect 34412 75124 34468 75518
rect 34412 75058 34468 75068
rect 34972 76636 35252 76692
rect 35644 77588 35700 77598
rect 34188 74900 34244 74910
rect 34524 74900 34580 74910
rect 34188 74898 34356 74900
rect 34188 74846 34190 74898
rect 34242 74846 34356 74898
rect 34188 74844 34356 74846
rect 34188 74834 34244 74844
rect 34076 74722 34132 74732
rect 34188 74340 34244 74350
rect 34188 74246 34244 74284
rect 33852 74162 33908 74172
rect 34300 74228 34356 74844
rect 33292 73892 33348 73902
rect 33292 73444 33348 73836
rect 33404 73892 33460 73902
rect 33404 73890 33908 73892
rect 33404 73838 33406 73890
rect 33458 73838 33908 73890
rect 33404 73836 33908 73838
rect 33404 73826 33460 73836
rect 33740 73668 33796 73678
rect 33628 73556 33684 73566
rect 33628 73462 33684 73500
rect 33404 73444 33460 73454
rect 33292 73388 33404 73444
rect 33068 72658 33348 72660
rect 33068 72606 33070 72658
rect 33122 72606 33348 72658
rect 33068 72604 33348 72606
rect 33068 72594 33124 72604
rect 33292 72436 33348 72604
rect 33404 72658 33460 73388
rect 33404 72606 33406 72658
rect 33458 72606 33460 72658
rect 33404 72594 33460 72606
rect 33740 72660 33796 73612
rect 33852 73330 33908 73836
rect 33852 73278 33854 73330
rect 33906 73278 33908 73330
rect 33852 73266 33908 73278
rect 33852 72660 33908 72670
rect 33740 72658 34020 72660
rect 33740 72606 33854 72658
rect 33906 72606 34020 72658
rect 33740 72604 34020 72606
rect 33852 72594 33908 72604
rect 33292 72380 33684 72436
rect 31948 72270 31950 72322
rect 32002 72270 32004 72322
rect 19836 72156 20100 72166
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 19836 72090 20100 72100
rect 4476 71372 4740 71382
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4476 71306 4740 71316
rect 19836 70588 20100 70598
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 19836 70522 20100 70532
rect 31948 70532 32004 72270
rect 33628 71202 33684 72380
rect 33964 71986 34020 72604
rect 33964 71934 33966 71986
rect 34018 71934 34020 71986
rect 33964 71922 34020 71934
rect 34300 71986 34356 74172
rect 34412 74844 34524 74900
rect 34412 73668 34468 74844
rect 34524 74806 34580 74844
rect 34636 74898 34692 74910
rect 34636 74846 34638 74898
rect 34690 74846 34692 74898
rect 34524 74228 34580 74238
rect 34524 74134 34580 74172
rect 34636 74004 34692 74846
rect 34636 73938 34692 73948
rect 34748 74116 34804 74126
rect 34412 73602 34468 73612
rect 34748 73556 34804 74060
rect 34860 73556 34916 73566
rect 34748 73554 34916 73556
rect 34748 73502 34862 73554
rect 34914 73502 34916 73554
rect 34748 73500 34916 73502
rect 34860 73490 34916 73500
rect 34524 73444 34580 73454
rect 34524 73350 34580 73388
rect 34972 72772 35028 76636
rect 35084 76466 35140 76478
rect 35084 76414 35086 76466
rect 35138 76414 35140 76466
rect 35084 75572 35140 76414
rect 35196 76076 35460 76086
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35196 76010 35460 76020
rect 35196 75572 35252 75582
rect 35532 75572 35588 75582
rect 35084 75570 35252 75572
rect 35084 75518 35198 75570
rect 35250 75518 35252 75570
rect 35084 75516 35252 75518
rect 35196 75506 35252 75516
rect 35308 75570 35588 75572
rect 35308 75518 35534 75570
rect 35586 75518 35588 75570
rect 35308 75516 35588 75518
rect 35308 75122 35364 75516
rect 35532 75506 35588 75516
rect 35644 75124 35700 77532
rect 35868 76354 35924 79200
rect 37212 76804 37268 79200
rect 37884 77026 37940 79200
rect 37884 76974 37886 77026
rect 37938 76974 37940 77026
rect 37884 76962 37940 76974
rect 35868 76302 35870 76354
rect 35922 76302 35924 76354
rect 35868 76290 35924 76302
rect 36988 76748 37268 76804
rect 36092 76020 36148 76030
rect 36092 75682 36148 75964
rect 36204 75908 36260 75918
rect 36204 75794 36260 75852
rect 36204 75742 36206 75794
rect 36258 75742 36260 75794
rect 36204 75730 36260 75742
rect 36092 75630 36094 75682
rect 36146 75630 36148 75682
rect 35308 75070 35310 75122
rect 35362 75070 35364 75122
rect 35308 75058 35364 75070
rect 35532 75068 35700 75124
rect 35756 75124 35812 75134
rect 36092 75124 36148 75630
rect 36764 75570 36820 75582
rect 36764 75518 36766 75570
rect 36818 75518 36820 75570
rect 36316 75458 36372 75470
rect 36316 75406 36318 75458
rect 36370 75406 36372 75458
rect 36316 75124 36372 75406
rect 36540 75460 36596 75470
rect 36540 75458 36708 75460
rect 36540 75406 36542 75458
rect 36594 75406 36708 75458
rect 36540 75404 36708 75406
rect 36540 75394 36596 75404
rect 36540 75124 36596 75134
rect 36092 75068 36260 75124
rect 36316 75122 36596 75124
rect 36316 75070 36542 75122
rect 36594 75070 36596 75122
rect 36316 75068 36596 75070
rect 35196 74508 35460 74518
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35196 74442 35460 74452
rect 35532 74340 35588 75068
rect 35308 74284 35588 74340
rect 35644 74900 35700 74910
rect 35644 74674 35700 74844
rect 35644 74622 35646 74674
rect 35698 74622 35700 74674
rect 35644 74452 35700 74622
rect 35308 74228 35364 74284
rect 35308 74114 35364 74172
rect 35308 74062 35310 74114
rect 35362 74062 35364 74114
rect 35308 74050 35364 74062
rect 35532 74116 35588 74126
rect 35644 74116 35700 74396
rect 35532 74114 35700 74116
rect 35532 74062 35534 74114
rect 35586 74062 35700 74114
rect 35532 74060 35700 74062
rect 35532 74050 35588 74060
rect 35420 74004 35476 74014
rect 35420 73910 35476 73948
rect 35756 73554 35812 75068
rect 36092 74900 36148 74910
rect 35868 74788 35924 74798
rect 35868 74786 36036 74788
rect 35868 74734 35870 74786
rect 35922 74734 36036 74786
rect 35868 74732 36036 74734
rect 35868 74722 35924 74732
rect 35980 74116 36036 74732
rect 35980 74022 36036 74060
rect 35756 73502 35758 73554
rect 35810 73502 35812 73554
rect 35756 73490 35812 73502
rect 35196 72940 35460 72950
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35196 72874 35460 72884
rect 34972 72716 35476 72772
rect 35084 72548 35140 72558
rect 35084 72454 35140 72492
rect 34412 72436 34468 72446
rect 34412 72342 34468 72380
rect 34524 72434 34580 72446
rect 34524 72382 34526 72434
rect 34578 72382 34580 72434
rect 34300 71934 34302 71986
rect 34354 71934 34356 71986
rect 33628 71150 33630 71202
rect 33682 71150 33684 71202
rect 33628 71138 33684 71150
rect 34300 71092 34356 71934
rect 34524 71876 34580 72382
rect 35196 72436 35252 72446
rect 35196 72342 35252 72380
rect 35420 71986 35476 72716
rect 35980 72436 36036 72446
rect 36092 72436 36148 74844
rect 36204 74004 36260 75068
rect 36540 75058 36596 75068
rect 36428 74788 36484 74798
rect 36204 73948 36372 74004
rect 35980 72434 36148 72436
rect 35980 72382 35982 72434
rect 36034 72382 36148 72434
rect 35980 72380 36148 72382
rect 36204 72660 36260 72670
rect 36204 72436 36260 72604
rect 35980 72370 36036 72380
rect 35420 71934 35422 71986
rect 35474 71934 35476 71986
rect 35420 71922 35476 71934
rect 36092 71988 36148 71998
rect 36204 71988 36260 72380
rect 36092 71986 36260 71988
rect 36092 71934 36094 71986
rect 36146 71934 36260 71986
rect 36092 71932 36260 71934
rect 36092 71922 36148 71932
rect 34748 71876 34804 71886
rect 34524 71820 34748 71876
rect 34748 71782 34804 71820
rect 35196 71372 35460 71382
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35196 71306 35460 71316
rect 34300 71026 34356 71036
rect 34748 71202 34804 71214
rect 34748 71150 34750 71202
rect 34802 71150 34804 71202
rect 34748 71090 34804 71150
rect 34748 71038 34750 71090
rect 34802 71038 34804 71090
rect 34748 71026 34804 71038
rect 35308 71092 35364 71102
rect 35308 70998 35364 71036
rect 31948 70466 32004 70476
rect 36316 70420 36372 73948
rect 36428 73554 36484 74732
rect 36540 74340 36596 74350
rect 36540 74114 36596 74284
rect 36540 74062 36542 74114
rect 36594 74062 36596 74114
rect 36540 74050 36596 74062
rect 36652 74116 36708 75404
rect 36764 74564 36820 75518
rect 36988 74900 37044 76748
rect 37212 76578 37268 76590
rect 38108 76580 38164 76590
rect 37212 76526 37214 76578
rect 37266 76526 37268 76578
rect 37100 76466 37156 76478
rect 37100 76414 37102 76466
rect 37154 76414 37156 76466
rect 37100 76356 37156 76414
rect 37212 76468 37268 76526
rect 37212 76402 37268 76412
rect 37996 76578 38164 76580
rect 37996 76526 38110 76578
rect 38162 76526 38164 76578
rect 37996 76524 38164 76526
rect 37100 76290 37156 76300
rect 37884 76356 37940 76366
rect 37884 76262 37940 76300
rect 37212 76244 37268 76254
rect 37212 76150 37268 76188
rect 37884 75908 37940 75918
rect 37996 75908 38052 76524
rect 38108 76514 38164 76524
rect 38556 76580 38612 79200
rect 37884 75906 38052 75908
rect 37884 75854 37886 75906
rect 37938 75854 38052 75906
rect 37884 75852 38052 75854
rect 38220 76242 38276 76254
rect 38220 76190 38222 76242
rect 38274 76190 38276 76242
rect 37884 75842 37940 75852
rect 38108 75684 38164 75694
rect 36988 74834 37044 74844
rect 37100 75682 38164 75684
rect 37100 75630 38110 75682
rect 38162 75630 38164 75682
rect 37100 75628 38164 75630
rect 36764 74498 36820 74508
rect 36876 74674 36932 74686
rect 36876 74622 36878 74674
rect 36930 74622 36932 74674
rect 36652 74060 36820 74116
rect 36428 73502 36430 73554
rect 36482 73502 36484 73554
rect 36428 73490 36484 73502
rect 36652 73890 36708 73902
rect 36652 73838 36654 73890
rect 36706 73838 36708 73890
rect 36652 73556 36708 73838
rect 36652 73490 36708 73500
rect 36764 73332 36820 74060
rect 36876 74114 36932 74622
rect 36876 74062 36878 74114
rect 36930 74062 36932 74114
rect 36876 74050 36932 74062
rect 36988 74564 37044 74574
rect 36540 73276 36820 73332
rect 36876 73892 36932 73902
rect 36540 72772 36596 73276
rect 36764 73106 36820 73118
rect 36764 73054 36766 73106
rect 36818 73054 36820 73106
rect 36540 72660 36596 72716
rect 36652 72772 36708 72782
rect 36764 72772 36820 73054
rect 36652 72770 36820 72772
rect 36652 72718 36654 72770
rect 36706 72718 36820 72770
rect 36652 72716 36820 72718
rect 36652 72706 36708 72716
rect 36428 72604 36596 72660
rect 36428 72324 36484 72604
rect 36876 72548 36932 73836
rect 36652 72492 36932 72548
rect 36540 72436 36596 72446
rect 36540 72342 36596 72380
rect 36652 72434 36708 72492
rect 36652 72382 36654 72434
rect 36706 72382 36708 72434
rect 36652 72370 36708 72382
rect 36428 72258 36484 72268
rect 36876 72324 36932 72334
rect 36428 72100 36484 72110
rect 36428 71986 36484 72044
rect 36428 71934 36430 71986
rect 36482 71934 36484 71986
rect 36428 71922 36484 71934
rect 36876 71316 36932 72268
rect 36988 71874 37044 74508
rect 37100 71986 37156 75628
rect 38108 75618 38164 75628
rect 37324 75460 37380 75470
rect 37100 71934 37102 71986
rect 37154 71934 37156 71986
rect 37100 71922 37156 71934
rect 37212 75458 37380 75460
rect 37212 75406 37326 75458
rect 37378 75406 37380 75458
rect 37212 75404 37380 75406
rect 36988 71822 36990 71874
rect 37042 71822 37044 71874
rect 36988 71810 37044 71822
rect 36428 71092 36484 71102
rect 36428 70998 36484 71036
rect 36876 71090 36932 71260
rect 36876 71038 36878 71090
rect 36930 71038 36932 71090
rect 36876 71026 36932 71038
rect 36316 70354 36372 70364
rect 37100 70420 37156 70430
rect 37100 70326 37156 70364
rect 37212 70196 37268 75404
rect 37324 75394 37380 75404
rect 37660 75460 37716 75470
rect 37660 75366 37716 75404
rect 37436 75012 37492 75022
rect 37324 75010 37492 75012
rect 37324 74958 37438 75010
rect 37490 74958 37492 75010
rect 37324 74956 37492 74958
rect 37324 71988 37380 74956
rect 37436 74946 37492 74956
rect 37660 74898 37716 74910
rect 37660 74846 37662 74898
rect 37714 74846 37716 74898
rect 37548 74116 37604 74126
rect 37548 74022 37604 74060
rect 37660 74116 37716 74846
rect 37884 74900 37940 74910
rect 37772 74116 37828 74126
rect 37660 74060 37772 74116
rect 37660 73892 37716 74060
rect 37772 74050 37828 74060
rect 37436 73836 37716 73892
rect 37436 73330 37492 73836
rect 37436 73278 37438 73330
rect 37490 73278 37492 73330
rect 37436 73266 37492 73278
rect 37548 73442 37604 73454
rect 37548 73390 37550 73442
rect 37602 73390 37604 73442
rect 37548 73332 37604 73390
rect 37548 73266 37604 73276
rect 37884 72996 37940 74844
rect 37996 74564 38052 74574
rect 37996 74226 38052 74508
rect 37996 74174 37998 74226
rect 38050 74174 38052 74226
rect 37996 74162 38052 74174
rect 38108 74116 38164 74126
rect 37996 74002 38052 74014
rect 37996 73950 37998 74002
rect 38050 73950 38052 74002
rect 37996 73780 38052 73950
rect 38108 74002 38164 74060
rect 38108 73950 38110 74002
rect 38162 73950 38164 74002
rect 38108 73938 38164 73950
rect 37996 73714 38052 73724
rect 38220 73668 38276 76190
rect 38444 74900 38500 74910
rect 38444 74806 38500 74844
rect 38556 74004 38612 76524
rect 38780 77026 38836 77038
rect 38780 76974 38782 77026
rect 38834 76974 38836 77026
rect 38780 75794 38836 76974
rect 38892 76580 38948 76590
rect 38892 76486 38948 76524
rect 39228 75908 39284 79200
rect 39564 76356 39620 76366
rect 39452 76244 39508 76254
rect 39228 75852 39396 75908
rect 38780 75742 38782 75794
rect 38834 75742 38836 75794
rect 38780 75730 38836 75742
rect 38780 75012 38836 75022
rect 38780 74918 38836 74956
rect 38892 74900 38948 74910
rect 38892 74114 38948 74844
rect 39340 74676 39396 75852
rect 39452 75796 39508 76188
rect 39452 75122 39508 75740
rect 39452 75070 39454 75122
rect 39506 75070 39508 75122
rect 39452 75058 39508 75070
rect 38892 74062 38894 74114
rect 38946 74062 38948 74114
rect 38892 74050 38948 74062
rect 39228 74620 39396 74676
rect 38444 73948 38612 74004
rect 39004 74004 39060 74042
rect 38220 73602 38276 73612
rect 38332 73890 38388 73902
rect 38332 73838 38334 73890
rect 38386 73838 38388 73890
rect 38220 73332 38276 73342
rect 38220 73238 38276 73276
rect 37772 72940 37940 72996
rect 37772 72546 37828 72940
rect 37772 72494 37774 72546
rect 37826 72494 37828 72546
rect 37436 72436 37492 72446
rect 37436 72342 37492 72380
rect 37660 72322 37716 72334
rect 37660 72270 37662 72322
rect 37714 72270 37716 72322
rect 37660 72212 37716 72270
rect 37660 72146 37716 72156
rect 37324 71922 37380 71932
rect 37548 72100 37604 72110
rect 37436 70308 37492 70318
rect 37436 70214 37492 70252
rect 37212 70130 37268 70140
rect 37548 69970 37604 72044
rect 37772 72100 37828 72494
rect 37772 72034 37828 72044
rect 37884 72436 37940 72446
rect 37772 71764 37828 71774
rect 37884 71764 37940 72380
rect 37996 72212 38052 72222
rect 37996 71986 38052 72156
rect 37996 71934 37998 71986
rect 38050 71934 38052 71986
rect 37996 71922 38052 71934
rect 38332 71988 38388 73838
rect 38332 71922 38388 71932
rect 37772 71762 37940 71764
rect 37772 71710 37774 71762
rect 37826 71710 37940 71762
rect 37772 71708 37940 71710
rect 37660 71092 37716 71102
rect 37772 71092 37828 71708
rect 37660 71090 37828 71092
rect 37660 71038 37662 71090
rect 37714 71038 37828 71090
rect 37660 71036 37828 71038
rect 37660 71026 37716 71036
rect 38108 70868 38164 70878
rect 38108 70774 38164 70812
rect 37996 70420 38052 70430
rect 38444 70420 38500 73948
rect 39004 73938 39060 73948
rect 39116 73890 39172 73902
rect 39116 73838 39118 73890
rect 39170 73838 39172 73890
rect 39116 73780 39172 73838
rect 38780 73724 39172 73780
rect 38668 73668 38724 73678
rect 38668 73332 38724 73612
rect 38668 73200 38724 73276
rect 38556 72212 38612 72222
rect 38556 71090 38612 72156
rect 38780 72212 38836 73724
rect 39228 73668 39284 74620
rect 39564 74114 39620 76300
rect 39788 75684 39844 75694
rect 39676 75348 39732 75358
rect 39676 75122 39732 75292
rect 39676 75070 39678 75122
rect 39730 75070 39732 75122
rect 39676 74900 39732 75070
rect 39788 75122 39844 75628
rect 39788 75070 39790 75122
rect 39842 75070 39844 75122
rect 39788 75058 39844 75070
rect 39900 75124 39956 79200
rect 40572 76580 40628 79200
rect 40572 76514 40628 76524
rect 41132 76580 41188 76590
rect 41244 76580 41300 79200
rect 41244 76524 41412 76580
rect 40124 76468 40180 76478
rect 40180 76412 40292 76468
rect 40124 76402 40180 76412
rect 40236 76356 40292 76412
rect 41020 76356 41076 76366
rect 40236 76354 40404 76356
rect 40236 76302 40238 76354
rect 40290 76302 40404 76354
rect 40236 76300 40404 76302
rect 40236 76290 40292 76300
rect 40348 76244 40404 76300
rect 41020 76262 41076 76300
rect 40348 76178 40404 76188
rect 40908 75908 40964 75918
rect 40460 75906 40964 75908
rect 40460 75854 40910 75906
rect 40962 75854 40964 75906
rect 40460 75852 40964 75854
rect 40012 75796 40068 75806
rect 40012 75570 40068 75740
rect 40460 75794 40516 75852
rect 40908 75842 40964 75852
rect 40460 75742 40462 75794
rect 40514 75742 40516 75794
rect 40460 75730 40516 75742
rect 40684 75684 40740 75694
rect 40684 75590 40740 75628
rect 40012 75518 40014 75570
rect 40066 75518 40068 75570
rect 40012 75506 40068 75518
rect 40796 75572 40852 75582
rect 40124 75458 40180 75470
rect 40124 75406 40126 75458
rect 40178 75406 40180 75458
rect 40124 75236 40180 75406
rect 40124 75170 40180 75180
rect 40236 75460 40292 75470
rect 39900 75058 39956 75068
rect 39676 74834 39732 74844
rect 39900 74900 39956 74910
rect 40236 74900 40292 75404
rect 40796 75122 40852 75516
rect 40796 75070 40798 75122
rect 40850 75070 40852 75122
rect 39900 74898 40292 74900
rect 39900 74846 39902 74898
rect 39954 74846 40292 74898
rect 39900 74844 40292 74846
rect 40460 75010 40516 75022
rect 40460 74958 40462 75010
rect 40514 74958 40516 75010
rect 39900 74834 39956 74844
rect 40124 74228 40180 74238
rect 40124 74134 40180 74172
rect 39564 74062 39566 74114
rect 39618 74062 39620 74114
rect 39564 73948 39620 74062
rect 40460 74116 40516 74958
rect 39564 73892 39732 73948
rect 39004 73612 39284 73668
rect 38892 72436 38948 72446
rect 38892 72342 38948 72380
rect 38780 72146 38836 72156
rect 38780 71762 38836 71774
rect 38780 71710 38782 71762
rect 38834 71710 38836 71762
rect 38780 71204 38836 71710
rect 38780 71138 38836 71148
rect 38556 71038 38558 71090
rect 38610 71038 38612 71090
rect 38556 70980 38612 71038
rect 38556 70914 38612 70924
rect 38780 70978 38836 70990
rect 38780 70926 38782 70978
rect 38834 70926 38836 70978
rect 38780 70868 38836 70926
rect 38780 70802 38836 70812
rect 37996 70418 38500 70420
rect 37996 70366 37998 70418
rect 38050 70366 38500 70418
rect 37996 70364 38500 70366
rect 39004 70418 39060 73612
rect 39116 73218 39172 73230
rect 39116 73166 39118 73218
rect 39170 73166 39172 73218
rect 39116 72772 39172 73166
rect 39116 72706 39172 72716
rect 39116 72546 39172 72558
rect 39116 72494 39118 72546
rect 39170 72494 39172 72546
rect 39116 71876 39172 72494
rect 39116 71820 39620 71876
rect 39116 71762 39172 71820
rect 39116 71710 39118 71762
rect 39170 71710 39172 71762
rect 39116 71698 39172 71710
rect 39228 71650 39284 71662
rect 39228 71598 39230 71650
rect 39282 71598 39284 71650
rect 39116 71204 39172 71214
rect 39228 71204 39284 71598
rect 39116 71202 39284 71204
rect 39116 71150 39118 71202
rect 39170 71150 39284 71202
rect 39116 71148 39284 71150
rect 39116 71138 39172 71148
rect 39004 70366 39006 70418
rect 39058 70366 39060 70418
rect 37996 70354 38052 70364
rect 39004 70354 39060 70366
rect 39564 70418 39620 71820
rect 39676 71428 39732 73892
rect 40236 73780 40292 73790
rect 40236 73554 40292 73724
rect 40236 73502 40238 73554
rect 40290 73502 40292 73554
rect 40236 73490 40292 73502
rect 40348 73556 40404 73566
rect 40460 73556 40516 74060
rect 40572 75012 40628 75022
rect 40572 74114 40628 74956
rect 40796 75012 40852 75070
rect 40796 74946 40852 74956
rect 40572 74062 40574 74114
rect 40626 74062 40628 74114
rect 40572 74004 40628 74062
rect 40572 73938 40628 73948
rect 40684 74340 40740 74350
rect 40684 74114 40740 74284
rect 40684 74062 40686 74114
rect 40738 74062 40740 74114
rect 40348 73554 40516 73556
rect 40348 73502 40350 73554
rect 40402 73502 40516 73554
rect 40348 73500 40516 73502
rect 40572 73556 40628 73566
rect 40348 73490 40404 73500
rect 40572 73462 40628 73500
rect 40684 73444 40740 74062
rect 40796 74116 40852 74126
rect 40796 74022 40852 74060
rect 41132 73948 41188 76524
rect 40908 73892 41188 73948
rect 41244 75458 41300 75470
rect 41244 75406 41246 75458
rect 41298 75406 41300 75458
rect 41244 74114 41300 75406
rect 41244 74062 41246 74114
rect 41298 74062 41300 74114
rect 40796 73444 40852 73454
rect 40684 73442 40852 73444
rect 40684 73390 40798 73442
rect 40850 73390 40852 73442
rect 40684 73388 40852 73390
rect 40796 73378 40852 73388
rect 40460 73332 40516 73342
rect 39788 73218 39844 73230
rect 39788 73166 39790 73218
rect 39842 73166 39844 73218
rect 39788 72548 39844 73166
rect 40236 72772 40292 72782
rect 40124 72548 40180 72558
rect 39788 72546 40180 72548
rect 39788 72494 40126 72546
rect 40178 72494 40180 72546
rect 39788 72492 40180 72494
rect 40124 71652 40180 72492
rect 40236 72322 40292 72716
rect 40236 72270 40238 72322
rect 40290 72270 40292 72322
rect 40236 72212 40292 72270
rect 40236 72156 40404 72212
rect 39676 71372 39844 71428
rect 39676 71204 39732 71214
rect 39676 71110 39732 71148
rect 39676 70980 39732 70990
rect 39676 70886 39732 70924
rect 39564 70366 39566 70418
rect 39618 70366 39620 70418
rect 39564 70354 39620 70366
rect 39676 70308 39732 70318
rect 39788 70308 39844 71372
rect 40012 71204 40068 71214
rect 40124 71204 40180 71596
rect 40348 71650 40404 72156
rect 40460 71762 40516 73276
rect 40460 71710 40462 71762
rect 40514 71710 40516 71762
rect 40460 71698 40516 71710
rect 40348 71598 40350 71650
rect 40402 71598 40404 71650
rect 40348 71586 40404 71598
rect 40012 71202 40180 71204
rect 40012 71150 40014 71202
rect 40066 71150 40180 71202
rect 40012 71148 40180 71150
rect 40236 71538 40292 71550
rect 40236 71486 40238 71538
rect 40290 71486 40292 71538
rect 40012 70868 40068 71148
rect 40236 71092 40292 71486
rect 40236 71026 40292 71036
rect 40012 70802 40068 70812
rect 40460 70868 40516 70878
rect 39676 70306 39844 70308
rect 39676 70254 39678 70306
rect 39730 70254 39844 70306
rect 39676 70252 39844 70254
rect 40348 70308 40404 70318
rect 39676 70242 39732 70252
rect 40348 70214 40404 70252
rect 40236 70196 40292 70206
rect 40236 70102 40292 70140
rect 37548 69918 37550 69970
rect 37602 69918 37604 69970
rect 37548 69906 37604 69918
rect 38332 70082 38388 70094
rect 38332 70030 38334 70082
rect 38386 70030 38388 70082
rect 38332 69970 38388 70030
rect 38332 69918 38334 69970
rect 38386 69918 38388 69970
rect 4476 69804 4740 69814
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4476 69738 4740 69748
rect 35196 69804 35460 69814
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35196 69738 35460 69748
rect 38332 69634 38388 69918
rect 38332 69582 38334 69634
rect 38386 69582 38388 69634
rect 38332 69570 38388 69582
rect 39788 69634 39844 69646
rect 39788 69582 39790 69634
rect 39842 69582 39844 69634
rect 39788 69522 39844 69582
rect 39788 69470 39790 69522
rect 39842 69470 39844 69522
rect 39788 69458 39844 69470
rect 40348 69524 40404 69534
rect 40460 69524 40516 70812
rect 40796 70308 40852 70318
rect 40796 70214 40852 70252
rect 40348 69522 40516 69524
rect 40348 69470 40350 69522
rect 40402 69470 40516 69522
rect 40348 69468 40516 69470
rect 40796 69524 40852 69534
rect 40908 69524 40964 73892
rect 41244 72212 41300 74062
rect 41244 72146 41300 72156
rect 41244 71764 41300 71774
rect 41020 71092 41076 71102
rect 41020 70998 41076 71036
rect 41244 70978 41300 71708
rect 41244 70926 41246 70978
rect 41298 70926 41300 70978
rect 41244 70914 41300 70926
rect 41356 70756 41412 76524
rect 41692 76468 41748 76478
rect 41468 76244 41524 76254
rect 41468 74900 41524 76188
rect 41692 76244 41748 76412
rect 41580 75906 41636 75918
rect 41580 75854 41582 75906
rect 41634 75854 41636 75906
rect 41580 75124 41636 75854
rect 41692 75348 41748 76188
rect 41804 75572 41860 75582
rect 41804 75478 41860 75516
rect 41692 75292 41860 75348
rect 41692 75124 41748 75134
rect 41580 75122 41748 75124
rect 41580 75070 41694 75122
rect 41746 75070 41748 75122
rect 41580 75068 41748 75070
rect 41692 75058 41748 75068
rect 41804 75122 41860 75292
rect 41804 75070 41806 75122
rect 41858 75070 41860 75122
rect 41804 75058 41860 75070
rect 41580 74900 41636 74910
rect 41468 74898 41636 74900
rect 41468 74846 41582 74898
rect 41634 74846 41636 74898
rect 41468 74844 41636 74846
rect 41580 74834 41636 74844
rect 41692 74900 41748 74910
rect 41916 74900 41972 79200
rect 42028 76580 42084 76590
rect 42028 76486 42084 76524
rect 42588 76580 42644 79200
rect 43260 76692 43316 79200
rect 42588 76514 42644 76524
rect 43148 76636 43316 76692
rect 43372 76692 43428 76702
rect 43036 76468 43092 76478
rect 43036 76374 43092 76412
rect 42476 76132 42532 76142
rect 42252 75572 42308 75582
rect 42140 75460 42196 75470
rect 42252 75460 42308 75516
rect 42140 75458 42308 75460
rect 42140 75406 42142 75458
rect 42194 75406 42308 75458
rect 42140 75404 42308 75406
rect 42140 75394 42196 75404
rect 41916 74844 42084 74900
rect 41580 74116 41636 74126
rect 41692 74116 41748 74844
rect 42028 74452 42084 74844
rect 41636 74060 41748 74116
rect 41580 74050 41636 74060
rect 41468 73556 41524 73566
rect 41468 73462 41524 73500
rect 41692 73554 41748 74060
rect 41916 74396 42084 74452
rect 42140 74452 42196 74462
rect 41692 73502 41694 73554
rect 41746 73502 41748 73554
rect 41692 73490 41748 73502
rect 41804 74004 41860 74014
rect 41804 73442 41860 73948
rect 41916 73780 41972 74396
rect 42140 74226 42196 74396
rect 42140 74174 42142 74226
rect 42194 74174 42196 74226
rect 42140 74162 42196 74174
rect 42252 74340 42308 75404
rect 41916 73714 41972 73724
rect 42028 74114 42084 74126
rect 42028 74062 42030 74114
rect 42082 74062 42084 74114
rect 41804 73390 41806 73442
rect 41858 73390 41860 73442
rect 41804 73378 41860 73390
rect 41804 72996 41860 73006
rect 41580 72548 41636 72558
rect 41580 72454 41636 72492
rect 41692 72434 41748 72446
rect 41692 72382 41694 72434
rect 41746 72382 41748 72434
rect 41468 72324 41524 72334
rect 41468 72230 41524 72268
rect 41692 72324 41748 72382
rect 41692 72258 41748 72268
rect 41804 72436 41860 72940
rect 41804 72100 41860 72380
rect 41468 72044 41860 72100
rect 41916 72212 41972 72222
rect 41468 71986 41524 72044
rect 41468 71934 41470 71986
rect 41522 71934 41524 71986
rect 41468 71922 41524 71934
rect 41916 71652 41972 72156
rect 41916 71586 41972 71596
rect 41804 70980 41860 70990
rect 42028 70980 42084 74062
rect 42252 74002 42308 74284
rect 42252 73950 42254 74002
rect 42306 73950 42308 74002
rect 42252 73938 42308 73950
rect 42364 74900 42420 74910
rect 42364 73444 42420 74844
rect 42364 73378 42420 73388
rect 42476 72660 42532 76076
rect 43036 75684 43092 75694
rect 43036 75590 43092 75628
rect 42812 75572 42868 75582
rect 42812 75478 42868 75516
rect 42924 75570 42980 75582
rect 42924 75518 42926 75570
rect 42978 75518 42980 75570
rect 42924 75124 42980 75518
rect 42924 75058 42980 75068
rect 42700 74900 42756 74910
rect 42588 74898 42756 74900
rect 42588 74846 42702 74898
rect 42754 74846 42756 74898
rect 42588 74844 42756 74846
rect 42588 74004 42644 74844
rect 42700 74834 42756 74844
rect 42924 74898 42980 74910
rect 43148 74900 43204 76636
rect 43372 76598 43428 76636
rect 43260 76466 43316 76478
rect 43260 76414 43262 76466
rect 43314 76414 43316 76466
rect 43260 76132 43316 76414
rect 43484 76466 43540 76478
rect 43484 76414 43486 76466
rect 43538 76414 43540 76466
rect 43260 76066 43316 76076
rect 43372 76356 43428 76366
rect 42924 74846 42926 74898
rect 42978 74846 42980 74898
rect 42812 74786 42868 74798
rect 42812 74734 42814 74786
rect 42866 74734 42868 74786
rect 42700 74228 42756 74238
rect 42812 74228 42868 74734
rect 42700 74226 42868 74228
rect 42700 74174 42702 74226
rect 42754 74174 42868 74226
rect 42700 74172 42868 74174
rect 42924 74228 42980 74846
rect 43036 74844 43204 74900
rect 43260 75460 43316 75470
rect 43036 74452 43092 74844
rect 43260 74674 43316 75404
rect 43260 74622 43262 74674
rect 43314 74622 43316 74674
rect 43260 74610 43316 74622
rect 43036 74396 43316 74452
rect 42700 74162 42756 74172
rect 42924 74162 42980 74172
rect 43036 74116 43092 74126
rect 43036 74022 43092 74060
rect 42700 74004 42756 74014
rect 42588 73948 42700 74004
rect 42476 72594 42532 72604
rect 42588 73218 42644 73230
rect 42588 73166 42590 73218
rect 42642 73166 42644 73218
rect 42588 72548 42644 73166
rect 42588 72482 42644 72492
rect 42700 72546 42756 73948
rect 43260 73668 43316 74396
rect 43260 73602 43316 73612
rect 43148 73220 43204 73230
rect 42812 73108 42868 73118
rect 42812 73014 42868 73052
rect 43036 73106 43092 73118
rect 43036 73054 43038 73106
rect 43090 73054 43092 73106
rect 42700 72494 42702 72546
rect 42754 72494 42756 72546
rect 42700 72482 42756 72494
rect 42252 72434 42308 72446
rect 42252 72382 42254 72434
rect 42306 72382 42308 72434
rect 41804 70978 42084 70980
rect 41804 70926 41806 70978
rect 41858 70926 42084 70978
rect 41804 70924 42084 70926
rect 42140 71762 42196 71774
rect 42140 71710 42142 71762
rect 42194 71710 42196 71762
rect 42140 71092 42196 71710
rect 42252 71764 42308 72382
rect 43036 72436 43092 73054
rect 43148 72658 43204 73164
rect 43148 72606 43150 72658
rect 43202 72606 43204 72658
rect 43148 72594 43204 72606
rect 43036 72370 43092 72380
rect 42252 71698 42308 71708
rect 42364 71988 42420 71998
rect 41804 70914 41860 70924
rect 41356 70700 41636 70756
rect 41580 70418 41636 70700
rect 41580 70366 41582 70418
rect 41634 70366 41636 70418
rect 41580 70354 41636 70366
rect 42140 70196 42196 71036
rect 42364 71090 42420 71932
rect 42364 71038 42366 71090
rect 42418 71038 42420 71090
rect 42364 71026 42420 71038
rect 42924 71764 42980 71774
rect 43036 71764 43092 71774
rect 42980 71762 43092 71764
rect 42980 71710 43038 71762
rect 43090 71710 43092 71762
rect 42980 71708 43092 71710
rect 42812 70978 42868 70990
rect 42812 70926 42814 70978
rect 42866 70926 42868 70978
rect 42700 70420 42756 70430
rect 42812 70420 42868 70926
rect 42700 70418 42868 70420
rect 42700 70366 42702 70418
rect 42754 70366 42868 70418
rect 42700 70364 42868 70366
rect 42700 70354 42756 70364
rect 42364 70196 42420 70206
rect 42140 70194 42420 70196
rect 42140 70142 42366 70194
rect 42418 70142 42420 70194
rect 42140 70140 42420 70142
rect 42364 70130 42420 70140
rect 42812 70196 42868 70206
rect 42924 70196 42980 71708
rect 43036 71698 43092 71708
rect 43372 70644 43428 76300
rect 43484 75906 43540 76414
rect 43484 75854 43486 75906
rect 43538 75854 43540 75906
rect 43484 75842 43540 75854
rect 43596 76466 43652 76478
rect 43596 76414 43598 76466
rect 43650 76414 43652 76466
rect 43596 75908 43652 76414
rect 43596 75842 43652 75852
rect 43596 75124 43652 75134
rect 43484 74898 43540 74910
rect 43484 74846 43486 74898
rect 43538 74846 43540 74898
rect 43484 73556 43540 74846
rect 43484 73490 43540 73500
rect 43596 73332 43652 75068
rect 43932 74676 43988 79200
rect 44604 76692 44660 79200
rect 45276 76804 45332 79200
rect 45164 76748 45332 76804
rect 45388 77026 45444 77038
rect 45388 76974 45390 77026
rect 45442 76974 45444 77026
rect 44604 76626 44660 76636
rect 45052 76692 45108 76702
rect 44940 76578 44996 76590
rect 44940 76526 44942 76578
rect 44994 76526 44996 76578
rect 44716 76468 44772 76478
rect 44268 76356 44324 76366
rect 44268 75796 44324 76300
rect 44268 75730 44324 75740
rect 44156 75684 44212 75694
rect 44044 75460 44100 75470
rect 44044 75366 44100 75404
rect 43932 74610 43988 74620
rect 44156 74898 44212 75628
rect 44380 75570 44436 75582
rect 44380 75518 44382 75570
rect 44434 75518 44436 75570
rect 44380 75236 44436 75518
rect 44380 75170 44436 75180
rect 44268 75124 44324 75134
rect 44268 75030 44324 75068
rect 44716 75124 44772 76412
rect 44716 75058 44772 75068
rect 44828 76244 44884 76254
rect 44156 74846 44158 74898
rect 44210 74846 44212 74898
rect 44044 74228 44100 74238
rect 44044 74134 44100 74172
rect 43932 74116 43988 74126
rect 43932 74022 43988 74060
rect 44156 73892 44212 74846
rect 44492 74900 44548 74910
rect 44380 74452 44436 74462
rect 44268 74340 44324 74350
rect 44268 74246 44324 74284
rect 44380 74338 44436 74396
rect 44380 74286 44382 74338
rect 44434 74286 44436 74338
rect 43932 73836 44212 73892
rect 44380 74004 44436 74286
rect 44492 74116 44548 74844
rect 44716 74898 44772 74910
rect 44716 74846 44718 74898
rect 44770 74846 44772 74898
rect 44716 74340 44772 74846
rect 44716 74274 44772 74284
rect 44492 74050 44548 74060
rect 43820 73556 43876 73566
rect 43484 73276 43652 73332
rect 43708 73500 43820 73556
rect 43484 73106 43540 73276
rect 43484 73054 43486 73106
rect 43538 73054 43540 73106
rect 43484 73042 43540 73054
rect 43596 73108 43652 73118
rect 43596 71988 43652 73052
rect 43596 71894 43652 71932
rect 43708 72100 43764 73500
rect 43820 73462 43876 73500
rect 43932 72658 43988 73836
rect 43932 72606 43934 72658
rect 43986 72606 43988 72658
rect 43932 72594 43988 72606
rect 44268 73220 44324 73230
rect 44044 72548 44100 72558
rect 44044 72454 44100 72492
rect 43372 70578 43428 70588
rect 43484 71874 43540 71886
rect 43484 71822 43486 71874
rect 43538 71822 43540 71874
rect 43484 70420 43540 71822
rect 43708 71764 43764 72044
rect 43820 72322 43876 72334
rect 43820 72270 43822 72322
rect 43874 72270 43876 72322
rect 43820 71988 43876 72270
rect 43820 71922 43876 71932
rect 44156 72324 44212 72334
rect 44156 71874 44212 72268
rect 44156 71822 44158 71874
rect 44210 71822 44212 71874
rect 43820 71764 43876 71774
rect 43708 71762 43876 71764
rect 43708 71710 43822 71762
rect 43874 71710 43876 71762
rect 43708 71708 43876 71710
rect 43820 71092 43876 71708
rect 43820 71026 43876 71036
rect 44156 71090 44212 71822
rect 44156 71038 44158 71090
rect 44210 71038 44212 71090
rect 44156 71026 44212 71038
rect 44268 70868 44324 73164
rect 43932 70812 44324 70868
rect 43596 70420 43652 70430
rect 43036 70418 43652 70420
rect 43036 70366 43598 70418
rect 43650 70366 43652 70418
rect 43036 70364 43652 70366
rect 43036 70306 43092 70364
rect 43596 70354 43652 70364
rect 43036 70254 43038 70306
rect 43090 70254 43092 70306
rect 43036 70242 43092 70254
rect 42812 70194 42980 70196
rect 42812 70142 42814 70194
rect 42866 70142 42980 70194
rect 42812 70140 42980 70142
rect 43932 70194 43988 70812
rect 43932 70142 43934 70194
rect 43986 70142 43988 70194
rect 42812 70130 42868 70140
rect 43932 70130 43988 70142
rect 44156 70196 44212 70206
rect 44380 70196 44436 73948
rect 44604 73892 44660 73902
rect 44604 73330 44660 73836
rect 44604 73278 44606 73330
rect 44658 73278 44660 73330
rect 44604 72996 44660 73278
rect 44604 72930 44660 72940
rect 44828 73106 44884 76188
rect 44940 74452 44996 76526
rect 44940 74386 44996 74396
rect 44828 73054 44830 73106
rect 44882 73054 44884 73106
rect 44492 72548 44548 72558
rect 44492 72454 44548 72492
rect 44492 71092 44548 71102
rect 44492 70978 44548 71036
rect 44492 70926 44494 70978
rect 44546 70926 44548 70978
rect 44492 70914 44548 70926
rect 44716 71092 44772 71102
rect 44716 70418 44772 71036
rect 44716 70366 44718 70418
rect 44770 70366 44772 70418
rect 44716 70354 44772 70366
rect 44828 70308 44884 73054
rect 44940 72548 44996 72558
rect 44940 71986 44996 72492
rect 44940 71934 44942 71986
rect 44994 71934 44996 71986
rect 44940 71922 44996 71934
rect 44940 71764 44996 71774
rect 45052 71764 45108 76636
rect 45164 75460 45220 76748
rect 45276 76580 45332 76590
rect 45276 76486 45332 76524
rect 45164 75394 45220 75404
rect 45388 73668 45444 76974
rect 45836 76578 45892 76590
rect 45836 76526 45838 76578
rect 45890 76526 45892 76578
rect 45836 76244 45892 76526
rect 45948 76356 46004 79200
rect 46620 77252 46676 79200
rect 47180 77476 47236 77486
rect 46620 77196 47012 77252
rect 46732 77026 46788 77038
rect 46732 76974 46734 77026
rect 46786 76974 46788 77026
rect 46732 76690 46788 76974
rect 46732 76638 46734 76690
rect 46786 76638 46788 76690
rect 46732 76626 46788 76638
rect 46844 76580 46900 76590
rect 46172 76468 46228 76478
rect 46172 76466 46788 76468
rect 46172 76414 46174 76466
rect 46226 76414 46788 76466
rect 46172 76412 46788 76414
rect 45948 76300 46116 76356
rect 45836 76178 45892 76188
rect 45836 75570 45892 75582
rect 45836 75518 45838 75570
rect 45890 75518 45892 75570
rect 45500 75458 45556 75470
rect 45500 75406 45502 75458
rect 45554 75406 45556 75458
rect 45500 75348 45556 75406
rect 45500 75282 45556 75292
rect 45836 75124 45892 75518
rect 45836 75058 45892 75068
rect 45500 75012 45556 75022
rect 45500 74340 45556 74956
rect 45724 74900 45780 74910
rect 45724 74898 46004 74900
rect 45724 74846 45726 74898
rect 45778 74846 46004 74898
rect 45724 74844 46004 74846
rect 45724 74834 45780 74844
rect 45500 74274 45556 74284
rect 45612 74786 45668 74798
rect 45612 74734 45614 74786
rect 45666 74734 45668 74786
rect 45276 73612 45444 73668
rect 45276 73556 45332 73612
rect 45276 73490 45332 73500
rect 45388 73444 45444 73454
rect 45276 73332 45332 73370
rect 45388 73350 45444 73388
rect 45276 73266 45332 73276
rect 45276 73106 45332 73118
rect 45276 73054 45278 73106
rect 45330 73054 45332 73106
rect 45276 72772 45332 73054
rect 45612 73108 45668 74734
rect 45724 74340 45780 74350
rect 45724 74246 45780 74284
rect 45948 74226 46004 74844
rect 45948 74174 45950 74226
rect 46002 74174 46004 74226
rect 45948 73556 46004 74174
rect 45948 73490 46004 73500
rect 45836 73444 45892 73454
rect 45612 73052 45780 73108
rect 45276 72716 45668 72772
rect 45164 71988 45220 71998
rect 45276 71988 45332 72716
rect 45612 72546 45668 72716
rect 45612 72494 45614 72546
rect 45666 72494 45668 72546
rect 45612 72482 45668 72494
rect 45500 72434 45556 72446
rect 45500 72382 45502 72434
rect 45554 72382 45556 72434
rect 45500 72324 45556 72382
rect 45500 72258 45556 72268
rect 45724 72212 45780 73052
rect 45836 72884 45892 73388
rect 45948 73220 46004 73230
rect 45948 73126 46004 73164
rect 46060 73108 46116 76300
rect 46172 74898 46228 76412
rect 46284 76244 46340 76254
rect 46284 75794 46340 76188
rect 46732 75906 46788 76412
rect 46732 75854 46734 75906
rect 46786 75854 46788 75906
rect 46732 75842 46788 75854
rect 46844 76356 46900 76524
rect 46284 75742 46286 75794
rect 46338 75742 46340 75794
rect 46284 75730 46340 75742
rect 46844 75684 46900 76300
rect 46620 75628 46900 75684
rect 46172 74846 46174 74898
rect 46226 74846 46228 74898
rect 46172 74114 46228 74846
rect 46508 74898 46564 74910
rect 46508 74846 46510 74898
rect 46562 74846 46564 74898
rect 46172 74062 46174 74114
rect 46226 74062 46228 74114
rect 46172 74050 46228 74062
rect 46396 74116 46452 74126
rect 46284 73890 46340 73902
rect 46284 73838 46286 73890
rect 46338 73838 46340 73890
rect 46284 73218 46340 73838
rect 46396 73892 46452 74060
rect 46396 73826 46452 73836
rect 46508 73444 46564 74846
rect 46620 74116 46676 75628
rect 46956 75572 47012 77196
rect 47068 76692 47124 76702
rect 47068 76598 47124 76636
rect 47068 75572 47124 75582
rect 46956 75516 47068 75572
rect 47068 75506 47124 75516
rect 46844 75236 46900 75246
rect 46732 75124 46788 75134
rect 46732 75030 46788 75068
rect 46844 75010 46900 75180
rect 46844 74958 46846 75010
rect 46898 74958 46900 75010
rect 46844 74946 46900 74958
rect 47180 75124 47236 77420
rect 46620 74060 46900 74116
rect 46508 73378 46564 73388
rect 46732 73892 46788 73902
rect 46396 73332 46452 73342
rect 46396 73238 46452 73276
rect 46284 73166 46286 73218
rect 46338 73166 46340 73218
rect 46284 73154 46340 73166
rect 46060 73052 46228 73108
rect 45836 72828 46116 72884
rect 45724 72146 45780 72156
rect 45948 72212 46004 72222
rect 45164 71986 45332 71988
rect 45164 71934 45166 71986
rect 45218 71934 45332 71986
rect 45164 71932 45332 71934
rect 45836 72100 45892 72110
rect 45164 71922 45220 71932
rect 45276 71764 45332 71774
rect 45724 71764 45780 71774
rect 45052 71708 45220 71764
rect 44940 70420 44996 71708
rect 45052 70420 45108 70430
rect 44940 70418 45108 70420
rect 44940 70366 45054 70418
rect 45106 70366 45108 70418
rect 44940 70364 45108 70366
rect 45052 70354 45108 70364
rect 44828 70242 44884 70252
rect 44156 70194 44436 70196
rect 44156 70142 44158 70194
rect 44210 70142 44436 70194
rect 44156 70140 44436 70142
rect 44156 70130 44212 70140
rect 40796 69522 40964 69524
rect 40796 69470 40798 69522
rect 40850 69470 40964 69522
rect 40796 69468 40964 69470
rect 45164 69524 45220 71708
rect 45276 71762 45780 71764
rect 45276 71710 45278 71762
rect 45330 71710 45726 71762
rect 45778 71710 45780 71762
rect 45276 71708 45780 71710
rect 45276 71698 45332 71708
rect 45724 71698 45780 71708
rect 45388 71092 45444 71102
rect 45836 71092 45892 72044
rect 45948 71986 46004 72156
rect 45948 71934 45950 71986
rect 46002 71934 46004 71986
rect 45948 71922 46004 71934
rect 46060 71874 46116 72828
rect 46172 72772 46228 73052
rect 46172 72716 46676 72772
rect 46172 72546 46228 72558
rect 46172 72494 46174 72546
rect 46226 72494 46228 72546
rect 46172 72212 46228 72494
rect 46172 72146 46228 72156
rect 46620 71986 46676 72716
rect 46620 71934 46622 71986
rect 46674 71934 46676 71986
rect 46620 71922 46676 71934
rect 46060 71822 46062 71874
rect 46114 71822 46116 71874
rect 46060 71810 46116 71822
rect 45948 71092 46004 71102
rect 45836 71036 45948 71092
rect 45388 70998 45444 71036
rect 45948 70960 46004 71036
rect 46732 71090 46788 73836
rect 46844 72212 46900 74060
rect 47068 73890 47124 73902
rect 47068 73838 47070 73890
rect 47122 73838 47124 73890
rect 47068 73780 47124 73838
rect 47068 73714 47124 73724
rect 47068 73556 47124 73566
rect 47068 72770 47124 73500
rect 47068 72718 47070 72770
rect 47122 72718 47124 72770
rect 47068 72706 47124 72718
rect 46844 72146 46900 72156
rect 47180 72658 47236 75068
rect 47292 73332 47348 79200
rect 47964 77252 48020 79200
rect 47964 77196 48356 77252
rect 48076 77026 48132 77038
rect 48076 76974 48078 77026
rect 48130 76974 48132 77026
rect 47740 76578 47796 76590
rect 47740 76526 47742 76578
rect 47794 76526 47796 76578
rect 47516 76020 47572 76030
rect 47516 75122 47572 75964
rect 47516 75070 47518 75122
rect 47570 75070 47572 75122
rect 47516 75058 47572 75070
rect 47516 74676 47572 74686
rect 47516 73554 47572 74620
rect 47740 74116 47796 76526
rect 48076 76578 48132 76974
rect 48076 76526 48078 76578
rect 48130 76526 48132 76578
rect 47852 76244 47908 76254
rect 47852 74898 47908 76188
rect 47852 74846 47854 74898
rect 47906 74846 47908 74898
rect 47852 74834 47908 74846
rect 47740 74050 47796 74060
rect 47852 74452 47908 74462
rect 47740 73890 47796 73902
rect 47740 73838 47742 73890
rect 47794 73838 47796 73890
rect 47740 73668 47796 73838
rect 47740 73602 47796 73612
rect 47516 73502 47518 73554
rect 47570 73502 47572 73554
rect 47516 73490 47572 73502
rect 47292 73276 47796 73332
rect 47180 72606 47182 72658
rect 47234 72606 47236 72658
rect 46732 71038 46734 71090
rect 46786 71038 46788 71090
rect 46284 70754 46340 70766
rect 46284 70702 46286 70754
rect 46338 70702 46340 70754
rect 45500 70532 45556 70542
rect 45500 70418 45556 70476
rect 45500 70366 45502 70418
rect 45554 70366 45556 70418
rect 45500 70354 45556 70366
rect 46284 70308 46340 70702
rect 46396 70532 46452 70542
rect 46396 70418 46452 70476
rect 46396 70366 46398 70418
rect 46450 70366 46452 70418
rect 46396 70354 46452 70366
rect 46732 70420 46788 71038
rect 47180 71092 47236 72606
rect 47740 72434 47796 73276
rect 47740 72382 47742 72434
rect 47794 72382 47796 72434
rect 47740 72370 47796 72382
rect 47292 72212 47348 72222
rect 47292 71986 47348 72156
rect 47292 71934 47294 71986
rect 47346 71934 47348 71986
rect 47292 71922 47348 71934
rect 47740 72212 47796 72222
rect 47740 71986 47796 72156
rect 47740 71934 47742 71986
rect 47794 71934 47796 71986
rect 47740 71922 47796 71934
rect 47404 71092 47460 71102
rect 47180 71090 47460 71092
rect 47180 71038 47406 71090
rect 47458 71038 47460 71090
rect 47180 71036 47460 71038
rect 46844 70420 46900 70430
rect 46732 70418 46900 70420
rect 46732 70366 46846 70418
rect 46898 70366 46900 70418
rect 46732 70364 46900 70366
rect 46844 70354 46900 70364
rect 47180 70418 47236 71036
rect 47404 71026 47460 71036
rect 47852 71090 47908 74396
rect 47852 71038 47854 71090
rect 47906 71038 47908 71090
rect 47852 70980 47908 71038
rect 47852 70532 47908 70924
rect 47852 70466 47908 70476
rect 47180 70366 47182 70418
rect 47234 70366 47236 70418
rect 46284 70242 46340 70252
rect 40348 69458 40404 69468
rect 40796 69458 40852 69468
rect 45164 69458 45220 69468
rect 46172 70196 46228 70206
rect 46172 69522 46228 70140
rect 47180 70196 47236 70366
rect 48076 70420 48132 76526
rect 48188 75572 48244 75582
rect 48188 71876 48244 75516
rect 48300 72436 48356 77196
rect 48636 77026 48692 79200
rect 48636 76974 48638 77026
rect 48690 76974 48692 77026
rect 48636 76962 48692 76974
rect 49308 77028 49364 79200
rect 49308 76962 49364 76972
rect 49980 76804 50036 79200
rect 50652 77140 50708 79200
rect 49308 76748 50036 76804
rect 50428 77084 50652 77140
rect 48972 76580 49028 76590
rect 48972 76486 49028 76524
rect 49084 76468 49140 76478
rect 49084 76374 49140 76412
rect 48972 76244 49028 76254
rect 48972 76150 49028 76188
rect 48860 75572 48916 75582
rect 48860 75478 48916 75516
rect 49084 75460 49140 75470
rect 48412 75236 48468 75246
rect 48412 74338 48468 75180
rect 48636 75012 48692 75022
rect 48636 74918 48692 74956
rect 48524 74900 48580 74910
rect 48524 74806 48580 74844
rect 48412 74286 48414 74338
rect 48466 74286 48468 74338
rect 48412 74274 48468 74286
rect 48524 74452 48580 74462
rect 48524 74226 48580 74396
rect 48524 74174 48526 74226
rect 48578 74174 48580 74226
rect 48524 74162 48580 74174
rect 49084 73890 49140 75404
rect 49084 73838 49086 73890
rect 49138 73838 49140 73890
rect 49084 73826 49140 73838
rect 49196 74900 49252 74910
rect 48524 73442 48580 73454
rect 48524 73390 48526 73442
rect 48578 73390 48580 73442
rect 48412 72436 48468 72446
rect 48300 72434 48468 72436
rect 48300 72382 48414 72434
rect 48466 72382 48468 72434
rect 48300 72380 48468 72382
rect 48412 72370 48468 72380
rect 48524 72324 48580 73390
rect 48748 73444 48804 73454
rect 48748 73350 48804 73388
rect 48636 73220 48692 73230
rect 48636 73126 48692 73164
rect 48524 72258 48580 72268
rect 48636 72436 48692 72446
rect 48636 71986 48692 72380
rect 48636 71934 48638 71986
rect 48690 71934 48692 71986
rect 48188 71820 48356 71876
rect 48188 71650 48244 71662
rect 48188 71598 48190 71650
rect 48242 71598 48244 71650
rect 48188 71538 48244 71598
rect 48188 71486 48190 71538
rect 48242 71486 48244 71538
rect 48188 71474 48244 71486
rect 48300 71090 48356 71820
rect 48636 71538 48692 71934
rect 48636 71486 48638 71538
rect 48690 71486 48692 71538
rect 48636 71474 48692 71486
rect 48300 71038 48302 71090
rect 48354 71038 48356 71090
rect 48300 71026 48356 71038
rect 49196 71202 49252 74844
rect 49308 72434 49364 76748
rect 49868 76580 49924 76590
rect 49868 76486 49924 76524
rect 50092 76578 50148 76590
rect 50092 76526 50094 76578
rect 50146 76526 50148 76578
rect 49644 76468 49700 76478
rect 49644 75796 49700 76412
rect 49980 76354 50036 76366
rect 49980 76302 49982 76354
rect 50034 76302 50036 76354
rect 49644 75730 49700 75740
rect 49756 76244 49812 76254
rect 49756 75794 49812 76188
rect 49756 75742 49758 75794
rect 49810 75742 49812 75794
rect 49756 75236 49812 75742
rect 49308 72382 49310 72434
rect 49362 72382 49364 72434
rect 49308 72370 49364 72382
rect 49420 75180 49812 75236
rect 49868 75908 49924 75918
rect 49420 73332 49476 75180
rect 49532 74898 49588 74910
rect 49532 74846 49534 74898
rect 49586 74846 49588 74898
rect 49532 74788 49588 74846
rect 49532 74228 49588 74732
rect 49756 74340 49812 74350
rect 49868 74340 49924 75852
rect 49980 75010 50036 76302
rect 49980 74958 49982 75010
rect 50034 74958 50036 75010
rect 49980 74946 50036 74958
rect 50092 75572 50148 76526
rect 50092 75122 50148 75516
rect 50092 75070 50094 75122
rect 50146 75070 50148 75122
rect 50092 74900 50148 75070
rect 50092 74834 50148 74844
rect 50316 75012 50372 75022
rect 50428 75012 50484 77084
rect 50652 77074 50708 77084
rect 50556 76860 50820 76870
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50556 76794 50820 76804
rect 50764 76580 50820 76590
rect 50764 76486 50820 76524
rect 50988 76578 51044 76590
rect 50988 76526 50990 76578
rect 51042 76526 51044 76578
rect 50988 76356 51044 76526
rect 50988 76290 51044 76300
rect 51100 76466 51156 76478
rect 51100 76414 51102 76466
rect 51154 76414 51156 76466
rect 50876 75796 50932 75806
rect 50876 75702 50932 75740
rect 50764 75684 50820 75694
rect 50764 75590 50820 75628
rect 50988 75684 51044 75694
rect 51100 75684 51156 76414
rect 50988 75682 51156 75684
rect 50988 75630 50990 75682
rect 51042 75630 51156 75682
rect 50988 75628 51156 75630
rect 50988 75618 51044 75628
rect 50540 75460 50596 75470
rect 50540 75458 50932 75460
rect 50540 75406 50542 75458
rect 50594 75406 50932 75458
rect 50540 75404 50932 75406
rect 50540 75394 50596 75404
rect 50876 75348 50932 75404
rect 50556 75292 50820 75302
rect 50876 75292 51044 75348
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50556 75226 50820 75236
rect 50428 74956 50932 75012
rect 49756 74338 49924 74340
rect 49756 74286 49758 74338
rect 49810 74286 49924 74338
rect 49756 74284 49924 74286
rect 49980 74786 50036 74798
rect 49980 74734 49982 74786
rect 50034 74734 50036 74786
rect 49756 74274 49812 74284
rect 49532 74162 49588 74172
rect 49980 73556 50036 74734
rect 50316 74340 50372 74956
rect 49420 72436 49476 73276
rect 49420 72370 49476 72380
rect 49532 73500 50036 73556
rect 50092 74284 50372 74340
rect 50764 74788 50820 74798
rect 49532 71316 49588 73500
rect 50092 73444 50148 74284
rect 50540 74228 50596 74238
rect 49756 73388 50148 73444
rect 50204 74116 50260 74126
rect 50540 74114 50596 74172
rect 50204 74002 50260 74060
rect 50204 73950 50206 74002
rect 50258 73950 50260 74002
rect 49644 73220 49700 73230
rect 49644 73126 49700 73164
rect 49756 71874 49812 73388
rect 49980 73220 50036 73230
rect 49868 73106 49924 73118
rect 49868 73054 49870 73106
rect 49922 73054 49924 73106
rect 49868 72996 49924 73054
rect 49868 72546 49924 72940
rect 49868 72494 49870 72546
rect 49922 72494 49924 72546
rect 49868 72482 49924 72494
rect 49980 72548 50036 73164
rect 50092 73108 50148 73118
rect 50092 73014 50148 73052
rect 50092 72548 50148 72558
rect 49980 72546 50148 72548
rect 49980 72494 50094 72546
rect 50146 72494 50148 72546
rect 49980 72492 50148 72494
rect 50092 72482 50148 72492
rect 49980 72324 50036 72334
rect 50204 72324 50260 73950
rect 50316 74004 50372 74080
rect 50540 74062 50542 74114
rect 50594 74062 50596 74114
rect 50540 74050 50596 74062
rect 50316 73780 50372 73948
rect 50764 73892 50820 74732
rect 50764 73826 50820 73836
rect 50316 73724 50484 73780
rect 50428 73556 50484 73724
rect 50556 73724 50820 73734
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50556 73658 50820 73668
rect 50540 73556 50596 73566
rect 50428 73554 50596 73556
rect 50428 73502 50542 73554
rect 50594 73502 50596 73554
rect 50428 73500 50596 73502
rect 50540 73490 50596 73500
rect 50428 73108 50484 73118
rect 50428 72546 50484 73052
rect 50428 72494 50430 72546
rect 50482 72494 50484 72546
rect 50428 72482 50484 72494
rect 50876 72548 50932 74956
rect 50988 74788 51044 75292
rect 51100 75012 51156 75628
rect 51100 74946 51156 74956
rect 50988 74722 51044 74732
rect 51212 74786 51268 74798
rect 51212 74734 51214 74786
rect 51266 74734 51268 74786
rect 51212 74564 51268 74734
rect 51324 74676 51380 79200
rect 51660 76692 51716 76702
rect 51996 76692 52052 79200
rect 51660 76598 51716 76636
rect 51884 76636 52052 76692
rect 51772 76356 51828 76366
rect 51436 75684 51492 75694
rect 51772 75684 51828 76300
rect 51492 75682 51828 75684
rect 51492 75630 51774 75682
rect 51826 75630 51828 75682
rect 51492 75628 51828 75630
rect 51436 74900 51492 75628
rect 51772 75618 51828 75628
rect 51548 75460 51604 75470
rect 51548 75366 51604 75404
rect 51660 75458 51716 75470
rect 51660 75406 51662 75458
rect 51714 75406 51716 75458
rect 51660 75236 51716 75406
rect 51660 75170 51716 75180
rect 51772 75124 51828 75134
rect 51660 74900 51716 74910
rect 51436 74898 51716 74900
rect 51436 74846 51662 74898
rect 51714 74846 51716 74898
rect 51436 74844 51716 74846
rect 51324 74620 51492 74676
rect 50988 74508 51268 74564
rect 50988 73444 51044 74508
rect 51212 74340 51268 74350
rect 51100 74116 51156 74126
rect 51100 74022 51156 74060
rect 50988 73378 51044 73388
rect 51100 73444 51156 73454
rect 51212 73444 51268 74284
rect 51324 74004 51380 74014
rect 51324 73910 51380 73948
rect 51100 73442 51268 73444
rect 51100 73390 51102 73442
rect 51154 73390 51268 73442
rect 51100 73388 51268 73390
rect 51100 73378 51156 73388
rect 50988 73108 51044 73118
rect 50988 73014 51044 73052
rect 50876 72492 51044 72548
rect 49980 72322 50260 72324
rect 49980 72270 49982 72322
rect 50034 72270 50260 72322
rect 49980 72268 50260 72270
rect 50876 72324 50932 72334
rect 49980 72258 50036 72268
rect 50876 72230 50932 72268
rect 50556 72156 50820 72166
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50556 72090 50820 72100
rect 49756 71822 49758 71874
rect 49810 71822 49812 71874
rect 49756 71810 49812 71822
rect 50316 71764 50372 71774
rect 50316 71670 50372 71708
rect 49532 71250 49588 71260
rect 49196 71150 49198 71202
rect 49250 71150 49252 71202
rect 49196 71090 49252 71150
rect 50316 71202 50372 71214
rect 50316 71150 50318 71202
rect 50370 71150 50372 71202
rect 49196 71038 49198 71090
rect 49250 71038 49252 71090
rect 49196 71026 49252 71038
rect 49756 71092 49812 71102
rect 49756 70998 49812 71036
rect 50316 71092 50372 71150
rect 50876 71092 50932 71102
rect 50316 71090 50484 71092
rect 50316 71038 50318 71090
rect 50370 71038 50484 71090
rect 50316 71036 50484 71038
rect 50316 71026 50372 71036
rect 48748 70980 48804 70990
rect 48748 70886 48804 70924
rect 48412 70420 48468 70430
rect 48076 70418 48468 70420
rect 48076 70366 48414 70418
rect 48466 70366 48468 70418
rect 48076 70364 48468 70366
rect 48412 70354 48468 70364
rect 50428 70418 50484 71036
rect 50876 70998 50932 71036
rect 50556 70588 50820 70598
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50556 70522 50820 70532
rect 50428 70366 50430 70418
rect 50482 70366 50484 70418
rect 50428 70354 50484 70366
rect 47180 70130 47236 70140
rect 46172 69470 46174 69522
rect 46226 69470 46228 69522
rect 46172 69458 46228 69470
rect 46620 69524 46676 69534
rect 46620 69430 46676 69468
rect 50988 69524 51044 72492
rect 51324 72324 51380 72334
rect 51324 71762 51380 72268
rect 51324 71710 51326 71762
rect 51378 71710 51380 71762
rect 51324 70532 51380 71710
rect 51436 70868 51492 74620
rect 51548 74116 51604 74844
rect 51660 74834 51716 74844
rect 51660 74340 51716 74350
rect 51772 74340 51828 75068
rect 51884 74788 51940 76636
rect 51996 76468 52052 76478
rect 52108 76468 52164 76478
rect 51996 76466 52108 76468
rect 51996 76414 51998 76466
rect 52050 76414 52108 76466
rect 51996 76412 52108 76414
rect 51996 76402 52052 76412
rect 51996 76132 52052 76142
rect 51996 75124 52052 76076
rect 52108 75908 52164 76412
rect 52668 76468 52724 79200
rect 52668 76402 52724 76412
rect 52780 77364 52836 77374
rect 52668 76244 52724 76254
rect 52668 76150 52724 76188
rect 52556 76132 52612 76142
rect 52108 75852 52388 75908
rect 51996 75058 52052 75068
rect 52220 75682 52276 75694
rect 52220 75630 52222 75682
rect 52274 75630 52276 75682
rect 51884 74732 52052 74788
rect 51660 74338 51828 74340
rect 51660 74286 51662 74338
rect 51714 74286 51828 74338
rect 51660 74284 51828 74286
rect 51884 74564 51940 74574
rect 51660 74274 51716 74284
rect 51548 74060 51716 74116
rect 51548 73892 51604 73902
rect 51548 73798 51604 73836
rect 51548 70868 51604 70878
rect 51436 70866 51604 70868
rect 51436 70814 51550 70866
rect 51602 70814 51604 70866
rect 51436 70812 51604 70814
rect 51548 70802 51604 70812
rect 51324 70418 51380 70476
rect 51324 70366 51326 70418
rect 51378 70366 51380 70418
rect 51324 70354 51380 70366
rect 51660 70420 51716 74060
rect 51772 74004 51828 74014
rect 51772 73910 51828 73948
rect 51772 73444 51828 73454
rect 51772 71650 51828 73388
rect 51884 73330 51940 74508
rect 51996 73892 52052 74732
rect 52108 74786 52164 74798
rect 52108 74734 52110 74786
rect 52162 74734 52164 74786
rect 52108 74116 52164 74734
rect 52220 74340 52276 75630
rect 52220 74274 52276 74284
rect 52220 74116 52276 74126
rect 52108 74114 52276 74116
rect 52108 74062 52222 74114
rect 52274 74062 52276 74114
rect 52108 74060 52276 74062
rect 52220 74050 52276 74060
rect 51996 73836 52276 73892
rect 51884 73278 51886 73330
rect 51938 73278 51940 73330
rect 51884 72324 51940 73278
rect 52108 73218 52164 73230
rect 52108 73166 52110 73218
rect 52162 73166 52164 73218
rect 52108 72996 52164 73166
rect 52108 72930 52164 72940
rect 52108 72548 52164 72558
rect 52108 72454 52164 72492
rect 51884 72258 51940 72268
rect 51772 71598 51774 71650
rect 51826 71598 51828 71650
rect 51772 71586 51828 71598
rect 52220 70866 52276 73836
rect 52220 70814 52222 70866
rect 52274 70814 52276 70866
rect 52220 70802 52276 70814
rect 52220 70532 52276 70542
rect 51772 70420 51828 70430
rect 51660 70364 51772 70420
rect 51772 70288 51828 70364
rect 52220 70418 52276 70476
rect 52220 70366 52222 70418
rect 52274 70366 52276 70418
rect 52220 70354 52276 70366
rect 50988 69458 51044 69468
rect 52332 69522 52388 75852
rect 52556 75794 52612 76076
rect 52556 75742 52558 75794
rect 52610 75742 52612 75794
rect 52556 75730 52612 75742
rect 52444 75460 52500 75470
rect 52444 74116 52500 75404
rect 52780 74452 52836 77308
rect 53228 75124 53284 75134
rect 53340 75124 53396 79200
rect 53676 75684 53732 75694
rect 53676 75570 53732 75628
rect 53676 75518 53678 75570
rect 53730 75518 53732 75570
rect 53676 75506 53732 75518
rect 54012 75572 54068 79200
rect 54236 77588 54292 77598
rect 54124 75796 54180 75806
rect 54124 75702 54180 75740
rect 54012 75506 54068 75516
rect 53788 75458 53844 75470
rect 53788 75406 53790 75458
rect 53842 75406 53844 75458
rect 53340 75068 53732 75124
rect 53004 75010 53060 75022
rect 53004 74958 53006 75010
rect 53058 74958 53060 75010
rect 53004 74900 53060 74958
rect 53004 74834 53060 74844
rect 53228 74898 53284 75068
rect 53228 74846 53230 74898
rect 53282 74846 53284 74898
rect 53228 74834 53284 74846
rect 53564 74900 53620 74910
rect 52780 74386 52836 74396
rect 52556 74116 52612 74126
rect 53452 74116 53508 74126
rect 52444 74060 52556 74116
rect 52556 74022 52612 74060
rect 52668 74114 53508 74116
rect 52668 74062 53454 74114
rect 53506 74062 53508 74114
rect 52668 74060 53508 74062
rect 52444 73892 52500 73902
rect 52444 73556 52500 73836
rect 52444 73490 52500 73500
rect 52444 73332 52500 73342
rect 52444 72658 52500 73276
rect 52444 72606 52446 72658
rect 52498 72606 52500 72658
rect 52444 71874 52500 72606
rect 52556 73330 52612 73342
rect 52556 73278 52558 73330
rect 52610 73278 52612 73330
rect 52556 72548 52612 73278
rect 52556 72482 52612 72492
rect 52668 72546 52724 74060
rect 53452 74050 53508 74060
rect 53564 74004 53620 74844
rect 53564 73910 53620 73948
rect 53116 73556 53172 73566
rect 52780 73444 52836 73454
rect 52780 73442 52948 73444
rect 52780 73390 52782 73442
rect 52834 73390 52948 73442
rect 52780 73388 52948 73390
rect 52780 73378 52836 73388
rect 52668 72494 52670 72546
rect 52722 72494 52724 72546
rect 52668 72482 52724 72494
rect 52780 72548 52836 72558
rect 52444 71822 52446 71874
rect 52498 71822 52500 71874
rect 52444 71810 52500 71822
rect 52780 71874 52836 72492
rect 52780 71822 52782 71874
rect 52834 71822 52836 71874
rect 52780 71810 52836 71822
rect 52892 71988 52948 73388
rect 52556 71764 52612 71774
rect 52556 71670 52612 71708
rect 52892 71762 52948 71932
rect 52892 71710 52894 71762
rect 52946 71710 52948 71762
rect 52892 71698 52948 71710
rect 52668 70420 52724 70430
rect 52668 70326 52724 70364
rect 53116 70418 53172 73500
rect 53564 73332 53620 73342
rect 53564 73238 53620 73276
rect 53452 72548 53508 72558
rect 53452 72454 53508 72492
rect 53564 70868 53620 70878
rect 53676 70868 53732 75068
rect 53564 70866 53732 70868
rect 53564 70814 53566 70866
rect 53618 70814 53732 70866
rect 53564 70812 53732 70814
rect 53564 70802 53620 70812
rect 53116 70366 53118 70418
rect 53170 70366 53172 70418
rect 53116 70354 53172 70366
rect 53564 70420 53620 70430
rect 53564 70326 53620 70364
rect 53788 70308 53844 75406
rect 53900 75458 53956 75470
rect 53900 75406 53902 75458
rect 53954 75406 53956 75458
rect 53900 75124 53956 75406
rect 54236 75348 54292 77532
rect 53900 75058 53956 75068
rect 54012 75292 54292 75348
rect 54348 75682 54404 75694
rect 54348 75630 54350 75682
rect 54402 75630 54404 75682
rect 53900 74898 53956 74910
rect 53900 74846 53902 74898
rect 53954 74846 53956 74898
rect 53900 73108 53956 74846
rect 54012 74226 54068 75292
rect 54348 75236 54404 75630
rect 54684 75684 54740 79200
rect 54796 77140 54852 77150
rect 54796 76578 54852 77084
rect 55356 76692 55412 79200
rect 55356 76626 55412 76636
rect 55804 77028 55860 77038
rect 55804 76690 55860 76972
rect 56028 77028 56084 79200
rect 56028 76962 56084 76972
rect 55804 76638 55806 76690
rect 55858 76638 55860 76690
rect 55804 76626 55860 76638
rect 54796 76526 54798 76578
rect 54850 76526 54852 76578
rect 54796 76514 54852 76526
rect 56700 76580 56756 79200
rect 57372 76804 57428 79200
rect 57372 76738 57428 76748
rect 57596 77700 57652 77710
rect 56700 76514 56756 76524
rect 56924 76356 56980 76366
rect 56812 76354 56980 76356
rect 56812 76302 56926 76354
rect 56978 76302 56980 76354
rect 56812 76300 56980 76302
rect 56364 75908 56420 75918
rect 56364 75794 56420 75852
rect 56364 75742 56366 75794
rect 56418 75742 56420 75794
rect 56364 75730 56420 75742
rect 55916 75684 55972 75694
rect 54684 75628 55076 75684
rect 55020 75572 55076 75628
rect 55020 75570 55188 75572
rect 55020 75518 55022 75570
rect 55074 75518 55188 75570
rect 55020 75516 55188 75518
rect 55020 75506 55076 75516
rect 54348 75170 54404 75180
rect 54236 75122 54292 75134
rect 54236 75070 54238 75122
rect 54290 75070 54292 75122
rect 54124 75012 54180 75022
rect 54124 74918 54180 74956
rect 54012 74174 54014 74226
rect 54066 74174 54068 74226
rect 54012 74162 54068 74174
rect 54236 74226 54292 75070
rect 54348 75012 54404 75022
rect 54348 74898 54404 74956
rect 54348 74846 54350 74898
rect 54402 74846 54404 74898
rect 54348 74834 54404 74846
rect 54572 74900 54628 74910
rect 54236 74174 54238 74226
rect 54290 74174 54292 74226
rect 54236 74162 54292 74174
rect 54460 74114 54516 74126
rect 54460 74062 54462 74114
rect 54514 74062 54516 74114
rect 54460 73442 54516 74062
rect 54460 73390 54462 73442
rect 54514 73390 54516 73442
rect 54460 73378 54516 73390
rect 54572 73330 54628 74844
rect 54684 74898 54740 74910
rect 54684 74846 54686 74898
rect 54738 74846 54740 74898
rect 54684 74340 54740 74846
rect 54684 74274 54740 74284
rect 54572 73278 54574 73330
rect 54626 73278 54628 73330
rect 53900 72546 53956 73052
rect 54460 73108 54516 73118
rect 53900 72494 53902 72546
rect 53954 72494 53956 72546
rect 53900 72482 53956 72494
rect 54348 72660 54404 72670
rect 53900 71988 53956 71998
rect 53900 71894 53956 71932
rect 54236 71764 54292 71774
rect 54348 71764 54404 72604
rect 54236 71762 54404 71764
rect 54236 71710 54238 71762
rect 54290 71710 54404 71762
rect 54236 71708 54404 71710
rect 54460 71762 54516 73052
rect 54572 72996 54628 73278
rect 54796 74004 54852 74014
rect 54796 73330 54852 73948
rect 54796 73278 54798 73330
rect 54850 73278 54852 73330
rect 54796 73266 54852 73278
rect 54908 73108 54964 73118
rect 54908 73014 54964 73052
rect 54572 72940 54852 72996
rect 54796 72772 54852 72940
rect 54796 72716 55076 72772
rect 55020 72434 55076 72716
rect 55020 72382 55022 72434
rect 55074 72382 55076 72434
rect 55020 72370 55076 72382
rect 55132 72212 55188 75516
rect 55356 75236 55412 75246
rect 55356 75122 55412 75180
rect 55356 75070 55358 75122
rect 55410 75070 55412 75122
rect 55356 75058 55412 75070
rect 55244 75012 55300 75022
rect 55244 74918 55300 74956
rect 55468 74900 55524 74910
rect 55468 74806 55524 74844
rect 55916 74898 55972 75628
rect 56140 75460 56196 75470
rect 55916 74846 55918 74898
rect 55970 74846 55972 74898
rect 55916 74834 55972 74846
rect 56028 74900 56084 74910
rect 55468 74116 55524 74126
rect 55468 74022 55524 74060
rect 55916 74114 55972 74126
rect 55916 74062 55918 74114
rect 55970 74062 55972 74114
rect 55468 73668 55524 73678
rect 55468 73554 55524 73612
rect 55468 73502 55470 73554
rect 55522 73502 55524 73554
rect 55468 73490 55524 73502
rect 55804 73108 55860 73118
rect 55804 72772 55860 73052
rect 55804 72658 55860 72716
rect 55804 72606 55806 72658
rect 55858 72606 55860 72658
rect 55804 72594 55860 72606
rect 55356 72548 55412 72558
rect 55356 72454 55412 72492
rect 54460 71710 54462 71762
rect 54514 71710 54516 71762
rect 54236 71698 54292 71708
rect 54460 71202 54516 71710
rect 54460 71150 54462 71202
rect 54514 71150 54516 71202
rect 54460 71138 54516 71150
rect 54572 72156 55188 72212
rect 55356 72212 55412 72222
rect 54124 70754 54180 70766
rect 54124 70702 54126 70754
rect 54178 70702 54180 70754
rect 54124 70532 54180 70702
rect 54124 70466 54180 70476
rect 54572 70418 54628 72156
rect 55244 71764 55300 71774
rect 55356 71764 55412 72156
rect 55916 72212 55972 74062
rect 56028 74004 56084 74844
rect 56140 74338 56196 75404
rect 56364 75012 56420 75022
rect 56364 74918 56420 74956
rect 56700 75012 56756 75022
rect 56700 74918 56756 74956
rect 56140 74286 56142 74338
rect 56194 74286 56196 74338
rect 56140 74274 56196 74286
rect 56364 74452 56420 74462
rect 56028 73330 56084 73948
rect 56364 74226 56420 74396
rect 56364 74174 56366 74226
rect 56418 74174 56420 74226
rect 56252 73892 56308 73902
rect 56140 73556 56196 73566
rect 56140 73462 56196 73500
rect 56252 73554 56308 73836
rect 56252 73502 56254 73554
rect 56306 73502 56308 73554
rect 56028 73278 56030 73330
rect 56082 73278 56084 73330
rect 56028 72548 56084 73278
rect 56028 72482 56084 72492
rect 55916 72146 55972 72156
rect 55244 71762 55412 71764
rect 55244 71710 55246 71762
rect 55298 71710 55412 71762
rect 55244 71708 55412 71710
rect 55468 71874 55524 71886
rect 55468 71822 55470 71874
rect 55522 71822 55524 71874
rect 55468 71764 55524 71822
rect 56028 71764 56084 71774
rect 56252 71764 56308 73502
rect 55468 71762 56308 71764
rect 55468 71710 56030 71762
rect 56082 71710 56308 71762
rect 55468 71708 56308 71710
rect 55244 71698 55300 71708
rect 54684 71202 54740 71214
rect 54684 71150 54686 71202
rect 54738 71150 54740 71202
rect 54684 71090 54740 71150
rect 54684 71038 54686 71090
rect 54738 71038 54740 71090
rect 54684 71026 54740 71038
rect 55020 71202 55076 71214
rect 55020 71150 55022 71202
rect 55074 71150 55076 71202
rect 54572 70366 54574 70418
rect 54626 70366 54628 70418
rect 54572 70354 54628 70366
rect 55020 70418 55076 71150
rect 55244 71202 55300 71214
rect 55244 71150 55246 71202
rect 55298 71150 55300 71202
rect 55244 71090 55300 71150
rect 55244 71038 55246 71090
rect 55298 71038 55300 71090
rect 55244 71026 55300 71038
rect 55356 70980 55412 71708
rect 56028 71698 56084 71708
rect 56252 71540 56308 71550
rect 56252 71446 56308 71484
rect 55692 71092 55748 71102
rect 55692 70998 55748 71036
rect 55356 70914 55412 70924
rect 55580 70420 55636 70430
rect 55020 70366 55022 70418
rect 55074 70366 55076 70418
rect 55020 70354 55076 70366
rect 55468 70418 55636 70420
rect 55468 70366 55582 70418
rect 55634 70366 55636 70418
rect 55468 70364 55636 70366
rect 53788 70242 53844 70252
rect 55468 70306 55524 70364
rect 55580 70354 55636 70364
rect 56364 70418 56420 74174
rect 56700 73332 56756 73342
rect 56812 73332 56868 76300
rect 56924 76290 56980 76300
rect 57260 75908 57316 75918
rect 57148 75852 57260 75908
rect 56924 75796 56980 75806
rect 56924 75702 56980 75740
rect 57036 75460 57092 75470
rect 57036 75366 57092 75404
rect 57148 75236 57204 75852
rect 57260 75814 57316 75852
rect 57036 75180 57204 75236
rect 57036 74338 57092 75180
rect 57596 75122 57652 77644
rect 57932 76580 57988 76590
rect 57932 76486 57988 76524
rect 57596 75070 57598 75122
rect 57650 75070 57652 75122
rect 57596 75058 57652 75070
rect 57820 75458 57876 75470
rect 57820 75406 57822 75458
rect 57874 75406 57876 75458
rect 57036 74286 57038 74338
rect 57090 74286 57092 74338
rect 57036 74274 57092 74286
rect 57260 74228 57316 74238
rect 57260 74002 57316 74172
rect 57372 74228 57428 74238
rect 57372 74226 57764 74228
rect 57372 74174 57374 74226
rect 57426 74174 57764 74226
rect 57372 74172 57764 74174
rect 57372 74162 57428 74172
rect 57260 73950 57262 74002
rect 57314 73950 57316 74002
rect 57260 73938 57316 73950
rect 57596 73892 57652 73902
rect 57596 73554 57652 73836
rect 57596 73502 57598 73554
rect 57650 73502 57652 73554
rect 57596 73490 57652 73502
rect 56700 73330 56868 73332
rect 56700 73278 56702 73330
rect 56754 73278 56868 73330
rect 56700 73276 56868 73278
rect 57148 73332 57204 73342
rect 56700 72996 56756 73276
rect 56700 72930 56756 72940
rect 57148 72770 57204 73276
rect 57148 72718 57150 72770
rect 57202 72718 57204 72770
rect 57148 72706 57204 72718
rect 57484 73106 57540 73118
rect 57484 73054 57486 73106
rect 57538 73054 57540 73106
rect 56588 72658 56644 72670
rect 56588 72606 56590 72658
rect 56642 72606 56644 72658
rect 56588 71986 56644 72606
rect 56588 71934 56590 71986
rect 56642 71934 56644 71986
rect 56588 71922 56644 71934
rect 57036 72548 57092 72558
rect 56924 71092 56980 71102
rect 56924 70866 56980 71036
rect 57036 70978 57092 72492
rect 57484 72546 57540 73054
rect 57708 72772 57764 74172
rect 57820 74004 57876 75406
rect 58044 75236 58100 79200
rect 58716 76580 58772 79200
rect 58940 76580 58996 76590
rect 58716 76514 58772 76524
rect 58828 76578 58996 76580
rect 58828 76526 58942 76578
rect 58994 76526 58996 76578
rect 58828 76524 58996 76526
rect 58156 75572 58212 75582
rect 58156 75570 58324 75572
rect 58156 75518 58158 75570
rect 58210 75518 58324 75570
rect 58156 75516 58324 75518
rect 58156 75506 58212 75516
rect 58268 75460 58324 75516
rect 58268 75404 58436 75460
rect 58044 75170 58100 75180
rect 58156 75348 58212 75358
rect 58156 75010 58212 75292
rect 58156 74958 58158 75010
rect 58210 74958 58212 75010
rect 58156 74946 58212 74958
rect 57932 74676 57988 74686
rect 57932 74582 57988 74620
rect 57932 74004 57988 74014
rect 57820 73948 57932 74004
rect 57932 73910 57988 73948
rect 58268 74004 58324 74014
rect 58268 73910 58324 73948
rect 58044 73892 58100 73902
rect 58044 73798 58100 73836
rect 57820 73444 57876 73454
rect 57820 73350 57876 73388
rect 58268 73444 58324 73454
rect 57708 72716 58100 72772
rect 57484 72494 57486 72546
rect 57538 72494 57540 72546
rect 57484 72482 57540 72494
rect 57820 72546 57876 72558
rect 57820 72494 57822 72546
rect 57874 72494 57876 72546
rect 57036 70926 57038 70978
rect 57090 70926 57092 70978
rect 57036 70914 57092 70926
rect 57820 71650 57876 72494
rect 58044 72546 58100 72716
rect 58044 72494 58046 72546
rect 58098 72494 58100 72546
rect 58044 71762 58100 72494
rect 58044 71710 58046 71762
rect 58098 71710 58100 71762
rect 58044 71698 58100 71710
rect 57820 71598 57822 71650
rect 57874 71598 57876 71650
rect 56924 70814 56926 70866
rect 56978 70814 56980 70866
rect 56924 70802 56980 70814
rect 57820 70756 57876 71598
rect 58268 71540 58324 73388
rect 58380 73332 58436 75404
rect 58716 75458 58772 75470
rect 58716 75406 58718 75458
rect 58770 75406 58772 75458
rect 58716 75348 58772 75406
rect 58716 75282 58772 75292
rect 58380 73266 58436 73276
rect 58716 75010 58772 75022
rect 58716 74958 58718 75010
rect 58770 74958 58772 75010
rect 58604 73218 58660 73230
rect 58604 73166 58606 73218
rect 58658 73166 58660 73218
rect 58604 72660 58660 73166
rect 58604 72594 58660 72604
rect 58604 71876 58660 71886
rect 58716 71876 58772 74958
rect 58828 72772 58884 76524
rect 58940 76514 58996 76524
rect 59276 76580 59332 76590
rect 59276 76486 59332 76524
rect 59276 75796 59332 75806
rect 59052 75458 59108 75470
rect 59052 75406 59054 75458
rect 59106 75406 59108 75458
rect 58828 72706 58884 72716
rect 58940 75348 58996 75358
rect 58940 71988 58996 75292
rect 59052 74564 59108 75406
rect 59052 73556 59108 74508
rect 59164 74116 59220 74126
rect 59276 74116 59332 75740
rect 59388 75684 59444 79200
rect 59724 76356 59780 76366
rect 59724 76262 59780 76300
rect 59948 75796 60004 75806
rect 59388 75628 59780 75684
rect 59612 75460 59668 75470
rect 59612 75366 59668 75404
rect 59388 74898 59444 74910
rect 59388 74846 59390 74898
rect 59442 74846 59444 74898
rect 59388 74564 59444 74846
rect 59612 74898 59668 74910
rect 59612 74846 59614 74898
rect 59666 74846 59668 74898
rect 59388 74498 59444 74508
rect 59500 74786 59556 74798
rect 59500 74734 59502 74786
rect 59554 74734 59556 74786
rect 59388 74116 59444 74126
rect 59276 74114 59444 74116
rect 59276 74062 59390 74114
rect 59442 74062 59444 74114
rect 59276 74060 59444 74062
rect 59164 74022 59220 74060
rect 59388 74050 59444 74060
rect 59276 73890 59332 73902
rect 59276 73838 59278 73890
rect 59330 73838 59332 73890
rect 59052 73500 59220 73556
rect 59052 73330 59108 73342
rect 59052 73278 59054 73330
rect 59106 73278 59108 73330
rect 59052 72660 59108 73278
rect 59052 72594 59108 72604
rect 59164 72324 59220 73500
rect 59276 73220 59332 73838
rect 59500 73444 59556 74734
rect 59500 73378 59556 73388
rect 59612 74114 59668 74846
rect 59612 74062 59614 74114
rect 59666 74062 59668 74114
rect 59388 73220 59444 73230
rect 59276 73218 59444 73220
rect 59276 73166 59390 73218
rect 59442 73166 59444 73218
rect 59276 73164 59444 73166
rect 59388 73154 59444 73164
rect 59388 72996 59444 73006
rect 59388 72658 59444 72940
rect 59612 72770 59668 74062
rect 59724 73892 59780 75628
rect 59948 75570 60004 75740
rect 59948 75518 59950 75570
rect 60002 75518 60004 75570
rect 59948 74898 60004 75518
rect 59948 74846 59950 74898
rect 60002 74846 60004 74898
rect 59948 74834 60004 74846
rect 59836 74564 59892 74574
rect 59836 74338 59892 74508
rect 59836 74286 59838 74338
rect 59890 74286 59892 74338
rect 59836 74274 59892 74286
rect 59724 73826 59780 73836
rect 59836 74116 59892 74126
rect 59612 72718 59614 72770
rect 59666 72718 59668 72770
rect 59612 72706 59668 72718
rect 59388 72606 59390 72658
rect 59442 72606 59444 72658
rect 59388 72594 59444 72606
rect 59836 72658 59892 74060
rect 60060 73780 60116 79200
rect 60732 77026 60788 79200
rect 60732 76974 60734 77026
rect 60786 76974 60788 77026
rect 60732 76962 60788 76974
rect 61292 77026 61348 77038
rect 61292 76974 61294 77026
rect 61346 76974 61348 77026
rect 61292 76692 61348 76974
rect 61180 76690 61348 76692
rect 61180 76638 61294 76690
rect 61346 76638 61348 76690
rect 61180 76636 61348 76638
rect 60956 76578 61012 76590
rect 60956 76526 60958 76578
rect 61010 76526 61012 76578
rect 60508 75572 60564 75582
rect 60508 75478 60564 75516
rect 60956 75348 61012 76526
rect 60508 75292 61012 75348
rect 60284 74676 60340 74686
rect 60284 74114 60340 74620
rect 60508 74116 60564 75292
rect 60620 75180 61012 75236
rect 60620 75122 60676 75180
rect 60620 75070 60622 75122
rect 60674 75070 60676 75122
rect 60620 75058 60676 75070
rect 60732 75012 60788 75022
rect 60732 74918 60788 74956
rect 60620 74676 60676 74686
rect 60620 74674 60788 74676
rect 60620 74622 60622 74674
rect 60674 74622 60788 74674
rect 60620 74620 60788 74622
rect 60620 74610 60676 74620
rect 60284 74062 60286 74114
rect 60338 74062 60340 74114
rect 60284 74050 60340 74062
rect 60396 74060 60564 74116
rect 60060 73714 60116 73724
rect 60284 73444 60340 73454
rect 60284 73350 60340 73388
rect 60396 73332 60452 74060
rect 60620 74004 60676 74014
rect 60620 73910 60676 73948
rect 60508 73890 60564 73902
rect 60508 73838 60510 73890
rect 60562 73838 60564 73890
rect 60508 73556 60564 73838
rect 60732 73668 60788 74620
rect 60732 73602 60788 73612
rect 60844 73780 60900 73790
rect 60508 73490 60564 73500
rect 60844 73554 60900 73724
rect 60844 73502 60846 73554
rect 60898 73502 60900 73554
rect 60844 73490 60900 73502
rect 60956 73556 61012 75180
rect 60956 73490 61012 73500
rect 61068 74564 61124 74574
rect 60396 73276 60564 73332
rect 60172 73106 60228 73118
rect 60172 73054 60174 73106
rect 60226 73054 60228 73106
rect 60172 72770 60228 73054
rect 60172 72718 60174 72770
rect 60226 72718 60228 72770
rect 60172 72706 60228 72718
rect 59836 72606 59838 72658
rect 59890 72606 59892 72658
rect 59276 72548 59332 72558
rect 59276 72454 59332 72492
rect 59164 72268 59668 72324
rect 59052 71988 59108 71998
rect 58940 71986 59108 71988
rect 58940 71934 59054 71986
rect 59106 71934 59108 71986
rect 58940 71932 59108 71934
rect 59052 71922 59108 71932
rect 59612 71986 59668 72268
rect 59612 71934 59614 71986
rect 59666 71934 59668 71986
rect 59612 71922 59668 71934
rect 58604 71874 58772 71876
rect 58604 71822 58606 71874
rect 58658 71822 58772 71874
rect 58604 71820 58772 71822
rect 58604 71810 58660 71820
rect 58268 70866 58324 71484
rect 58940 71092 58996 71102
rect 58940 70998 58996 71036
rect 59836 71092 59892 72606
rect 60284 72660 60340 72670
rect 60284 72566 60340 72604
rect 59836 71026 59892 71036
rect 58268 70814 58270 70866
rect 58322 70814 58324 70866
rect 58268 70802 58324 70814
rect 58156 70756 58212 70766
rect 57820 70754 58212 70756
rect 57820 70702 58158 70754
rect 58210 70702 58212 70754
rect 57820 70700 58212 70702
rect 58156 70690 58212 70700
rect 60508 70532 60564 73276
rect 61068 72660 61124 74508
rect 61180 74340 61236 76636
rect 61292 76626 61348 76636
rect 61292 75684 61348 75694
rect 61292 75590 61348 75628
rect 61404 75124 61460 79200
rect 61852 76692 61908 76702
rect 61852 76598 61908 76636
rect 61852 76244 61908 76254
rect 61628 75908 61684 75918
rect 61628 75682 61684 75852
rect 61628 75630 61630 75682
rect 61682 75630 61684 75682
rect 61628 75618 61684 75630
rect 61404 75058 61460 75068
rect 61516 75460 61572 75470
rect 61404 74900 61460 74910
rect 61516 74900 61572 75404
rect 61404 74898 61572 74900
rect 61404 74846 61406 74898
rect 61458 74846 61572 74898
rect 61404 74844 61572 74846
rect 61404 74834 61460 74844
rect 61180 74274 61236 74284
rect 61292 74674 61348 74686
rect 61292 74622 61294 74674
rect 61346 74622 61348 74674
rect 61292 74228 61348 74622
rect 61852 74452 61908 76188
rect 62076 75572 62132 79200
rect 62524 77028 62580 77038
rect 62524 76690 62580 76972
rect 62524 76638 62526 76690
rect 62578 76638 62580 76690
rect 62524 76626 62580 76638
rect 62076 75506 62132 75516
rect 62188 75682 62244 75694
rect 62188 75630 62190 75682
rect 62242 75630 62244 75682
rect 61964 75236 62020 75246
rect 61964 75122 62020 75180
rect 61964 75070 61966 75122
rect 62018 75070 62020 75122
rect 61964 75058 62020 75070
rect 62188 75012 62244 75630
rect 62412 75684 62468 75694
rect 62188 74946 62244 74956
rect 62300 75570 62356 75582
rect 62300 75518 62302 75570
rect 62354 75518 62356 75570
rect 62300 74676 62356 75518
rect 62300 74610 62356 74620
rect 61852 74228 61908 74396
rect 61964 74228 62020 74238
rect 61852 74226 62020 74228
rect 61852 74174 61966 74226
rect 62018 74174 62020 74226
rect 61852 74172 62020 74174
rect 61292 74162 61348 74172
rect 61852 74004 61908 74014
rect 61404 73892 61460 73902
rect 61404 73798 61460 73836
rect 61404 73556 61460 73566
rect 61404 73462 61460 73500
rect 61852 73554 61908 73948
rect 61852 73502 61854 73554
rect 61906 73502 61908 73554
rect 61852 73490 61908 73502
rect 61292 72660 61348 72670
rect 61068 72658 61348 72660
rect 61068 72606 61294 72658
rect 61346 72606 61348 72658
rect 61068 72604 61348 72606
rect 61292 72594 61348 72604
rect 61964 72660 62020 74172
rect 62412 74226 62468 75628
rect 62748 75348 62804 79200
rect 63196 76804 63252 76814
rect 63196 76690 63252 76748
rect 63196 76638 63198 76690
rect 63250 76638 63252 76690
rect 63196 76626 63252 76638
rect 62860 75796 62916 75806
rect 62860 75702 62916 75740
rect 62636 75124 62692 75134
rect 62636 75030 62692 75068
rect 62412 74174 62414 74226
rect 62466 74174 62468 74226
rect 62300 73556 62356 73566
rect 62412 73556 62468 74174
rect 62356 73500 62468 73556
rect 62748 73556 62804 75292
rect 63308 75572 63364 75582
rect 63308 75122 63364 75516
rect 63308 75070 63310 75122
rect 63362 75070 63364 75122
rect 63308 75058 63364 75070
rect 63420 75124 63476 79200
rect 63756 76468 63812 76478
rect 63756 76374 63812 76412
rect 64092 75460 64148 79200
rect 64428 76580 64484 76590
rect 64428 76486 64484 76524
rect 64764 76580 64820 79200
rect 64764 75796 64820 76524
rect 64764 75730 64820 75740
rect 64876 76242 64932 76254
rect 64876 76190 64878 76242
rect 64930 76190 64932 76242
rect 64092 75394 64148 75404
rect 63420 75058 63476 75068
rect 63980 75124 64036 75134
rect 63980 75030 64036 75068
rect 64540 74786 64596 74798
rect 64540 74734 64542 74786
rect 64594 74734 64596 74786
rect 62860 74676 62916 74686
rect 62860 74226 62916 74620
rect 64540 74676 64596 74734
rect 64540 74610 64596 74620
rect 62860 74174 62862 74226
rect 62914 74174 62916 74226
rect 62860 74162 62916 74174
rect 63308 74340 63364 74350
rect 63308 74226 63364 74284
rect 63308 74174 63310 74226
rect 63362 74174 63364 74226
rect 63308 74162 63364 74174
rect 64876 74004 64932 76190
rect 65324 75796 65380 75806
rect 64988 75570 65044 75582
rect 64988 75518 64990 75570
rect 65042 75518 65044 75570
rect 64988 75348 65044 75518
rect 64988 75282 65044 75292
rect 65324 75124 65380 75740
rect 65436 75572 65492 79200
rect 66108 76244 66164 79200
rect 66108 76188 66388 76244
rect 65916 76076 66180 76086
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 65916 76010 66180 76020
rect 65436 75506 65492 75516
rect 65996 75460 66052 75470
rect 65996 75366 66052 75404
rect 66332 75460 66388 76188
rect 66780 75796 66836 79200
rect 67228 76580 67284 76590
rect 67228 76486 67284 76524
rect 66780 75730 66836 75740
rect 66668 75572 66724 75582
rect 66668 75478 66724 75516
rect 67452 75572 67508 79200
rect 67452 75506 67508 75516
rect 68012 75572 68068 75582
rect 68012 75478 68068 75516
rect 66332 75394 66388 75404
rect 67340 75460 67396 75470
rect 68124 75460 68180 79200
rect 68348 76244 68404 76254
rect 68348 76150 68404 76188
rect 68684 75796 68740 75806
rect 68684 75702 68740 75740
rect 68796 75460 68852 79200
rect 69356 76356 69412 76366
rect 69356 75570 69412 76300
rect 69356 75518 69358 75570
rect 69410 75518 69412 75570
rect 69356 75506 69412 75518
rect 69468 75572 69524 79200
rect 70140 76580 70196 79200
rect 70140 76514 70196 76524
rect 70588 76578 70644 76590
rect 70588 76526 70590 76578
rect 70642 76526 70644 76578
rect 70588 75796 70644 76526
rect 70588 75730 70644 75740
rect 69468 75506 69524 75516
rect 70252 75572 70308 75582
rect 70252 75478 70308 75516
rect 70812 75572 70868 79200
rect 70924 77476 70980 77486
rect 70924 75906 70980 77420
rect 71484 76804 71540 79200
rect 72156 76916 72212 79200
rect 72156 76850 72212 76860
rect 71484 76738 71540 76748
rect 72380 76804 72436 76814
rect 72380 76690 72436 76748
rect 72380 76638 72382 76690
rect 72434 76638 72436 76690
rect 72380 76626 72436 76638
rect 71484 76580 71540 76590
rect 71484 76486 71540 76524
rect 72828 76468 72884 79200
rect 73052 77364 73108 77374
rect 73052 76690 73108 77308
rect 73052 76638 73054 76690
rect 73106 76638 73108 76690
rect 73052 76626 73108 76638
rect 73500 76692 73556 79200
rect 74172 77250 74228 79200
rect 74172 77198 74174 77250
rect 74226 77198 74228 77250
rect 74172 77186 74228 77198
rect 73500 76626 73556 76636
rect 73948 76916 74004 76926
rect 73948 76690 74004 76860
rect 73948 76638 73950 76690
rect 74002 76638 74004 76690
rect 73948 76626 74004 76638
rect 74620 76692 74676 76702
rect 74620 76598 74676 76636
rect 73276 76468 73332 76478
rect 72828 76466 73332 76468
rect 72828 76414 73278 76466
rect 73330 76414 73332 76466
rect 72828 76412 73332 76414
rect 70924 75854 70926 75906
rect 70978 75854 70980 75906
rect 70924 75842 70980 75854
rect 68124 75404 68404 75460
rect 67340 75366 67396 75404
rect 65436 75124 65492 75134
rect 65324 75122 65492 75124
rect 65324 75070 65438 75122
rect 65490 75070 65492 75122
rect 65324 75068 65492 75070
rect 65436 75058 65492 75068
rect 68348 75122 68404 75404
rect 68796 75394 68852 75404
rect 69132 75460 69188 75470
rect 68348 75070 68350 75122
rect 68402 75070 68404 75122
rect 68348 75058 68404 75070
rect 69132 75122 69188 75404
rect 69692 75460 69748 75470
rect 69692 75366 69748 75404
rect 69132 75070 69134 75122
rect 69186 75070 69188 75122
rect 69132 75058 69188 75070
rect 70812 75122 70868 75516
rect 73052 75572 73108 75582
rect 73052 75478 73108 75516
rect 70812 75070 70814 75122
rect 70866 75070 70868 75122
rect 70812 75058 70868 75070
rect 73276 75122 73332 76412
rect 73948 75684 74004 75694
rect 73948 75590 74004 75628
rect 74844 75572 74900 79200
rect 75292 77250 75348 77262
rect 75292 77198 75294 77250
rect 75346 77198 75348 77250
rect 75292 76690 75348 77198
rect 75292 76638 75294 76690
rect 75346 76638 75348 76690
rect 75292 76626 75348 76638
rect 75516 76692 75572 79200
rect 76188 77026 76244 79200
rect 76188 76974 76190 77026
rect 76242 76974 76244 77026
rect 76188 76962 76244 76974
rect 75516 76626 75572 76636
rect 76300 76692 76356 76702
rect 76300 76598 76356 76636
rect 74844 75506 74900 75516
rect 76076 75572 76132 75582
rect 76076 75478 76132 75516
rect 73276 75070 73278 75122
rect 73330 75070 73332 75122
rect 73276 75058 73332 75070
rect 76860 75012 76916 79200
rect 76972 77026 77028 77038
rect 76972 76974 76974 77026
rect 77026 76974 77028 77026
rect 76972 76690 77028 76974
rect 76972 76638 76974 76690
rect 77026 76638 77028 76690
rect 76972 76626 77028 76638
rect 77532 76692 77588 79200
rect 77756 76692 77812 76702
rect 77532 76690 77812 76692
rect 77532 76638 77758 76690
rect 77810 76638 77812 76690
rect 77532 76636 77812 76638
rect 77756 76626 77812 76636
rect 77196 75572 77252 75582
rect 77196 75478 77252 75516
rect 78092 75572 78148 75582
rect 78204 75572 78260 79200
rect 78092 75570 78260 75572
rect 78092 75518 78094 75570
rect 78146 75518 78260 75570
rect 78092 75516 78260 75518
rect 78092 75506 78148 75516
rect 76860 74946 76916 74956
rect 77644 75012 77700 75022
rect 77644 74918 77700 74956
rect 78092 75012 78148 75022
rect 74508 74676 74564 74686
rect 74508 74582 74564 74620
rect 65916 74508 66180 74518
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 65916 74442 66180 74452
rect 78092 74226 78148 74956
rect 78092 74174 78094 74226
rect 78146 74174 78148 74226
rect 78092 74162 78148 74174
rect 64876 73938 64932 73948
rect 62860 73556 62916 73566
rect 62748 73554 62916 73556
rect 62748 73502 62862 73554
rect 62914 73502 62916 73554
rect 62748 73500 62916 73502
rect 62300 73424 62356 73500
rect 62860 73490 62916 73500
rect 65916 72940 66180 72950
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 65916 72874 66180 72884
rect 61964 72594 62020 72604
rect 65916 71372 66180 71382
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 65916 71306 66180 71316
rect 60508 70466 60564 70476
rect 56364 70366 56366 70418
rect 56418 70366 56420 70418
rect 56364 70354 56420 70366
rect 55468 70254 55470 70306
rect 55522 70254 55524 70306
rect 55468 70242 55524 70254
rect 65916 69804 66180 69814
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 65916 69738 66180 69748
rect 52332 69470 52334 69522
rect 52386 69470 52388 69522
rect 52332 69458 52388 69470
rect 52780 69524 52836 69534
rect 52780 69430 52836 69468
rect 19836 69020 20100 69030
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 19836 68954 20100 68964
rect 50556 69020 50820 69030
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50556 68954 50820 68964
rect 4476 68236 4740 68246
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4476 68170 4740 68180
rect 35196 68236 35460 68246
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35196 68170 35460 68180
rect 65916 68236 66180 68246
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 65916 68170 66180 68180
rect 19836 67452 20100 67462
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 19836 67386 20100 67396
rect 50556 67452 50820 67462
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50556 67386 50820 67396
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 35196 66668 35460 66678
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35196 66602 35460 66612
rect 65916 66668 66180 66678
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 65916 66602 66180 66612
rect 19836 65884 20100 65894
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 19836 65818 20100 65828
rect 50556 65884 50820 65894
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50556 65818 50820 65828
rect 4476 65100 4740 65110
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 35196 65100 35460 65110
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35196 65034 35460 65044
rect 65916 65100 66180 65110
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 65916 65034 66180 65044
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 50556 64316 50820 64326
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50556 64250 50820 64260
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35196 63466 35460 63476
rect 65916 63532 66180 63542
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 65916 63466 66180 63476
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 50556 62748 50820 62758
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50556 62682 50820 62692
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 65916 61964 66180 61974
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 65916 61898 66180 61908
rect 19836 61180 20100 61190
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 50556 61180 50820 61190
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50556 61114 50820 61124
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 65916 60396 66180 60406
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 65916 60330 66180 60340
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 50556 59612 50820 59622
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50556 59546 50820 59556
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 65916 58828 66180 58838
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 65916 58762 66180 58772
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 50556 58044 50820 58054
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50556 57978 50820 57988
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 65916 57260 66180 57270
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 65916 57194 66180 57204
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 65916 55692 66180 55702
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 65916 55626 66180 55636
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 65916 54124 66180 54134
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 65916 54058 66180 54068
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 65916 52556 66180 52566
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 65916 52490 66180 52500
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 65916 50988 66180 50998
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 65916 50922 66180 50932
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 65916 49420 66180 49430
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 65916 49354 66180 49364
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 65916 47852 66180 47862
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 65916 47786 66180 47796
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 65916 46284 66180 46294
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 65916 46218 66180 46228
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 65916 44716 66180 44726
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 65916 44650 66180 44660
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 65916 43148 66180 43158
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 65916 43082 66180 43092
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 65916 41580 66180 41590
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 65916 41514 66180 41524
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 65916 40012 66180 40022
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 65916 39946 66180 39956
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 65916 38444 66180 38454
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 65916 38378 66180 38388
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 65916 36876 66180 36886
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 65916 36810 66180 36820
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 65916 35308 66180 35318
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 65916 35242 66180 35252
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 65916 33740 66180 33750
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 65916 33674 66180 33684
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 65916 32172 66180 32182
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 65916 32106 66180 32116
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 65916 30604 66180 30614
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 65916 30538 66180 30548
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 65916 29036 66180 29046
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 65916 28970 66180 28980
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 65916 27468 66180 27478
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 65916 27402 66180 27412
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 65916 25900 66180 25910
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 65916 25834 66180 25844
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 65916 24332 66180 24342
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 65916 24266 66180 24276
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 65916 22764 66180 22774
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 65916 22698 66180 22708
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 65916 21196 66180 21206
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 65916 21130 66180 21140
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 65916 19628 66180 19638
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 65916 19562 66180 19572
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 65916 18060 66180 18070
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 65916 17994 66180 18004
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 65916 16492 66180 16502
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 65916 16426 66180 16436
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 65916 14924 66180 14934
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 65916 14858 66180 14868
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 65916 13356 66180 13366
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 65916 13290 66180 13300
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 65916 11788 66180 11798
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 65916 11722 66180 11732
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 65916 10220 66180 10230
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 65916 10154 66180 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 65916 8652 66180 8662
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 65916 8586 66180 8596
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 65916 7084 66180 7094
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 65916 7018 66180 7028
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 65916 5516 66180 5526
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 65916 5450 66180 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 13916 4452 13972 4462
rect 17948 4452 18004 4462
rect 24668 4452 24724 4462
rect 29372 4452 29428 4462
rect 32508 4452 32564 4462
rect 37212 4452 37268 4462
rect 51324 4452 51380 4462
rect 55356 4452 55412 4462
rect 59388 4452 59444 4462
rect 63420 4452 63476 4462
rect 70812 4452 70868 4462
rect 73388 4452 73444 4462
rect 13692 4450 13972 4452
rect 13692 4398 13918 4450
rect 13970 4398 13972 4450
rect 13692 4396 13972 4398
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 6972 3332 7028 3342
rect 6748 3330 7028 3332
rect 6748 3278 6974 3330
rect 7026 3278 7028 3330
rect 6748 3276 7028 3278
rect 6748 800 6804 3276
rect 6972 3266 7028 3276
rect 8092 3330 8148 3342
rect 8092 3278 8094 3330
rect 8146 3278 8148 3330
rect 8092 800 8148 3278
rect 8876 3332 8932 3342
rect 9996 3332 10052 3342
rect 8876 3330 9044 3332
rect 8876 3278 8878 3330
rect 8930 3278 9044 3330
rect 8876 3276 9044 3278
rect 8876 3266 8932 3276
rect 8988 800 9044 3276
rect 9884 3330 10052 3332
rect 9884 3278 9998 3330
rect 10050 3278 10052 3330
rect 9884 3276 10052 3278
rect 9884 800 9940 3276
rect 9996 3266 10052 3276
rect 10780 3330 10836 3342
rect 10780 3278 10782 3330
rect 10834 3278 10836 3330
rect 10780 800 10836 3278
rect 11452 3332 11508 3342
rect 12124 3332 12180 3342
rect 12796 3332 12852 3342
rect 11452 3330 11732 3332
rect 11452 3278 11454 3330
rect 11506 3278 11732 3330
rect 11452 3276 11732 3278
rect 11452 3266 11508 3276
rect 11676 800 11732 3276
rect 12124 3330 12404 3332
rect 12124 3278 12126 3330
rect 12178 3278 12404 3330
rect 12124 3276 12404 3278
rect 12124 3266 12180 3276
rect 12348 800 12404 3276
rect 12796 3330 13076 3332
rect 12796 3278 12798 3330
rect 12850 3278 13076 3330
rect 12796 3276 13076 3278
rect 12796 3266 12852 3276
rect 13020 800 13076 3276
rect 13692 800 13748 4396
rect 13916 4386 13972 4396
rect 17724 4450 18004 4452
rect 17724 4398 17950 4450
rect 18002 4398 18004 4450
rect 17724 4396 18004 4398
rect 14028 3332 14084 3342
rect 14700 3332 14756 3342
rect 15372 3332 15428 3342
rect 16044 3332 16100 3342
rect 16716 3332 16772 3342
rect 14028 3330 14420 3332
rect 14028 3278 14030 3330
rect 14082 3278 14420 3330
rect 14028 3276 14420 3278
rect 14028 3266 14084 3276
rect 14364 800 14420 3276
rect 14700 3330 15092 3332
rect 14700 3278 14702 3330
rect 14754 3278 15092 3330
rect 14700 3276 15092 3278
rect 14700 3266 14756 3276
rect 15036 800 15092 3276
rect 15372 3330 15764 3332
rect 15372 3278 15374 3330
rect 15426 3278 15764 3330
rect 15372 3276 15764 3278
rect 15372 3266 15428 3276
rect 15708 800 15764 3276
rect 16044 3330 16436 3332
rect 16044 3278 16046 3330
rect 16098 3278 16436 3330
rect 16044 3276 16436 3278
rect 16044 3266 16100 3276
rect 16380 800 16436 3276
rect 16716 3330 17108 3332
rect 16716 3278 16718 3330
rect 16770 3278 17108 3330
rect 16716 3276 17108 3278
rect 16716 3266 16772 3276
rect 17052 800 17108 3276
rect 17724 800 17780 4396
rect 17948 4386 18004 4396
rect 24444 4450 24724 4452
rect 24444 4398 24670 4450
rect 24722 4398 24724 4450
rect 24444 4396 24724 4398
rect 17948 3332 18004 3342
rect 18620 3332 18676 3342
rect 17948 3330 18452 3332
rect 17948 3278 17950 3330
rect 18002 3278 18452 3330
rect 17948 3276 18452 3278
rect 17948 3266 18004 3276
rect 18396 800 18452 3276
rect 18620 3330 19124 3332
rect 18620 3278 18622 3330
rect 18674 3278 19124 3330
rect 18620 3276 19124 3278
rect 18620 3266 18676 3276
rect 19068 800 19124 3276
rect 19292 3330 19348 3342
rect 19292 3278 19294 3330
rect 19346 3278 19348 3330
rect 19292 980 19348 3278
rect 19964 3332 20020 3342
rect 20636 3332 20692 3342
rect 19964 3330 20468 3332
rect 19964 3278 19966 3330
rect 20018 3278 20468 3330
rect 19964 3276 20468 3278
rect 19964 3266 20020 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 19292 924 19796 980
rect 19740 800 19796 924
rect 20412 800 20468 3276
rect 20636 3330 21140 3332
rect 20636 3278 20638 3330
rect 20690 3278 21140 3330
rect 20636 3276 21140 3278
rect 20636 3266 20692 3276
rect 21084 800 21140 3276
rect 21756 3330 21812 3342
rect 21756 3278 21758 3330
rect 21810 3278 21812 3330
rect 21756 800 21812 3278
rect 22428 3330 22484 3342
rect 22428 3278 22430 3330
rect 22482 3278 22484 3330
rect 22428 800 22484 3278
rect 23100 3330 23156 3342
rect 23100 3278 23102 3330
rect 23154 3278 23156 3330
rect 23100 800 23156 3278
rect 23772 3330 23828 3342
rect 23772 3278 23774 3330
rect 23826 3278 23828 3330
rect 23772 800 23828 3278
rect 24444 800 24500 4396
rect 24668 4386 24724 4396
rect 29148 4450 29428 4452
rect 29148 4398 29374 4450
rect 29426 4398 29428 4450
rect 29148 4396 29428 4398
rect 24556 3330 24612 3342
rect 24556 3278 24558 3330
rect 24610 3278 24612 3330
rect 24556 1762 24612 3278
rect 25788 3330 25844 3342
rect 25788 3278 25790 3330
rect 25842 3278 25844 3330
rect 24556 1710 24558 1762
rect 24610 1710 24612 1762
rect 24556 1698 24612 1710
rect 25116 1762 25172 1774
rect 25116 1710 25118 1762
rect 25170 1710 25172 1762
rect 25116 800 25172 1710
rect 25788 800 25844 3278
rect 26460 3330 26516 3342
rect 26460 3278 26462 3330
rect 26514 3278 26516 3330
rect 26460 800 26516 3278
rect 27132 3330 27188 3342
rect 27132 3278 27134 3330
rect 27186 3278 27188 3330
rect 27132 800 27188 3278
rect 27804 3330 27860 3342
rect 27804 3278 27806 3330
rect 27858 3278 27860 3330
rect 27804 800 27860 3278
rect 28476 3330 28532 3342
rect 28476 3278 28478 3330
rect 28530 3278 28532 3330
rect 28476 800 28532 3278
rect 29148 800 29204 4396
rect 29372 4386 29428 4396
rect 32284 4450 32564 4452
rect 32284 4398 32510 4450
rect 32562 4398 32564 4450
rect 32284 4396 32564 4398
rect 29708 3332 29764 3342
rect 29708 3330 29876 3332
rect 29708 3278 29710 3330
rect 29762 3278 29876 3330
rect 29708 3276 29876 3278
rect 29708 3266 29764 3276
rect 29820 800 29876 3276
rect 30268 3330 30324 3342
rect 30268 3278 30270 3330
rect 30322 3278 30324 3330
rect 30268 800 30324 3278
rect 30940 3330 30996 3342
rect 30940 3278 30942 3330
rect 30994 3278 30996 3330
rect 30940 800 30996 3278
rect 31612 3330 31668 3342
rect 31612 3278 31614 3330
rect 31666 3278 31668 3330
rect 31612 800 31668 3278
rect 32284 800 32340 4396
rect 32508 4386 32564 4396
rect 36988 4450 37268 4452
rect 36988 4398 37214 4450
rect 37266 4398 37268 4450
rect 36988 4396 37268 4398
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 32396 3330 32452 3342
rect 32396 3278 32398 3330
rect 32450 3278 32452 3330
rect 32396 1762 32452 3278
rect 33628 3330 33684 3342
rect 33628 3278 33630 3330
rect 33682 3278 33684 3330
rect 32396 1710 32398 1762
rect 32450 1710 32452 1762
rect 32396 1698 32452 1710
rect 32956 1762 33012 1774
rect 32956 1710 32958 1762
rect 33010 1710 33012 1762
rect 32956 800 33012 1710
rect 33628 800 33684 3278
rect 34300 3330 34356 3342
rect 34300 3278 34302 3330
rect 34354 3278 34356 3330
rect 34300 800 34356 3278
rect 34972 3330 35028 3342
rect 34972 3278 34974 3330
rect 35026 3278 35028 3330
rect 34972 800 35028 3278
rect 35644 3330 35700 3342
rect 35644 3278 35646 3330
rect 35698 3278 35700 3330
rect 35644 800 35700 3278
rect 36316 3330 36372 3342
rect 36316 3278 36318 3330
rect 36370 3278 36372 3330
rect 36316 800 36372 3278
rect 36988 800 37044 4396
rect 37212 4386 37268 4396
rect 51100 4450 51380 4452
rect 51100 4398 51326 4450
rect 51378 4398 51380 4450
rect 51100 4396 51380 4398
rect 37548 3332 37604 3342
rect 38220 3332 38276 3342
rect 38892 3332 38948 3342
rect 39564 3332 39620 3342
rect 40236 3332 40292 3342
rect 41244 3332 41300 3342
rect 41916 3332 41972 3342
rect 42588 3332 42644 3342
rect 43260 3332 43316 3342
rect 43932 3332 43988 3342
rect 37548 3330 37716 3332
rect 37548 3278 37550 3330
rect 37602 3278 37716 3330
rect 37548 3276 37716 3278
rect 37548 3266 37604 3276
rect 37660 800 37716 3276
rect 38220 3330 38388 3332
rect 38220 3278 38222 3330
rect 38274 3278 38388 3330
rect 38220 3276 38388 3278
rect 38220 3266 38276 3276
rect 38332 800 38388 3276
rect 38892 3330 39060 3332
rect 38892 3278 38894 3330
rect 38946 3278 39060 3330
rect 38892 3276 39060 3278
rect 38892 3266 38948 3276
rect 39004 800 39060 3276
rect 39564 3330 39732 3332
rect 39564 3278 39566 3330
rect 39618 3278 39732 3330
rect 39564 3276 39732 3278
rect 39564 3266 39620 3276
rect 39676 800 39732 3276
rect 40236 3330 40404 3332
rect 40236 3278 40238 3330
rect 40290 3278 40404 3330
rect 40236 3276 40404 3278
rect 40236 3266 40292 3276
rect 40348 800 40404 3276
rect 41020 3330 41300 3332
rect 41020 3278 41246 3330
rect 41298 3278 41300 3330
rect 41020 3276 41300 3278
rect 41020 800 41076 3276
rect 41244 3266 41300 3276
rect 41692 3330 41972 3332
rect 41692 3278 41918 3330
rect 41970 3278 41972 3330
rect 41692 3276 41972 3278
rect 41692 800 41748 3276
rect 41916 3266 41972 3276
rect 42364 3330 42644 3332
rect 42364 3278 42590 3330
rect 42642 3278 42644 3330
rect 42364 3276 42644 3278
rect 42364 800 42420 3276
rect 42588 3266 42644 3276
rect 43036 3330 43316 3332
rect 43036 3278 43262 3330
rect 43314 3278 43316 3330
rect 43036 3276 43316 3278
rect 43036 800 43092 3276
rect 43260 3266 43316 3276
rect 43708 3330 43988 3332
rect 43708 3278 43934 3330
rect 43986 3278 43988 3330
rect 43708 3276 43988 3278
rect 43708 800 43764 3276
rect 43932 3266 43988 3276
rect 44940 3330 44996 3342
rect 44940 3278 44942 3330
rect 44994 3278 44996 3330
rect 44380 1762 44436 1774
rect 44380 1710 44382 1762
rect 44434 1710 44436 1762
rect 44380 800 44436 1710
rect 44940 1762 44996 3278
rect 44940 1710 44942 1762
rect 44994 1710 44996 1762
rect 44940 1698 44996 1710
rect 45052 3332 45108 3342
rect 45052 800 45108 3276
rect 45612 3332 45668 3342
rect 45612 3238 45668 3276
rect 46284 3330 46340 3342
rect 46284 3278 46286 3330
rect 46338 3278 46340 3330
rect 45724 1762 45780 1774
rect 45724 1710 45726 1762
rect 45778 1710 45780 1762
rect 45724 800 45780 1710
rect 46284 1762 46340 3278
rect 46956 3330 47012 3342
rect 46956 3278 46958 3330
rect 47010 3278 47012 3330
rect 46284 1710 46286 1762
rect 46338 1710 46340 1762
rect 46284 1698 46340 1710
rect 46396 1874 46452 1886
rect 46396 1822 46398 1874
rect 46450 1822 46452 1874
rect 46396 800 46452 1822
rect 46956 1874 47012 3278
rect 46956 1822 46958 1874
rect 47010 1822 47012 1874
rect 46956 1810 47012 1822
rect 47628 3330 47684 3342
rect 47628 3278 47630 3330
rect 47682 3278 47684 3330
rect 47068 1762 47124 1774
rect 47068 1710 47070 1762
rect 47122 1710 47124 1762
rect 47068 800 47124 1710
rect 47628 1762 47684 3278
rect 47628 1710 47630 1762
rect 47682 1710 47684 1762
rect 47628 1698 47684 1710
rect 47740 3332 47796 3342
rect 47740 800 47796 3276
rect 48860 3332 48916 3342
rect 48860 3238 48916 3276
rect 49532 3330 49588 3342
rect 49532 3278 49534 3330
rect 49586 3278 49588 3330
rect 48412 1764 48468 1774
rect 48412 800 48468 1708
rect 49084 1762 49140 1774
rect 49084 1710 49086 1762
rect 49138 1710 49140 1762
rect 49084 800 49140 1710
rect 49532 1764 49588 3278
rect 49532 1698 49588 1708
rect 49756 3332 49812 3342
rect 49756 800 49812 3276
rect 50204 3330 50260 3342
rect 50204 3278 50206 3330
rect 50258 3278 50260 3330
rect 50204 1762 50260 3278
rect 50876 3332 50932 3342
rect 50876 3238 50932 3276
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 50204 1710 50206 1762
rect 50258 1710 50260 1762
rect 50204 1698 50260 1710
rect 50428 1762 50484 1774
rect 50428 1710 50430 1762
rect 50482 1710 50484 1762
rect 50428 800 50484 1710
rect 51100 800 51156 4396
rect 51324 4386 51380 4396
rect 55132 4450 55412 4452
rect 55132 4398 55358 4450
rect 55410 4398 55412 4450
rect 55132 4396 55412 4398
rect 51548 3330 51604 3342
rect 51548 3278 51550 3330
rect 51602 3278 51604 3330
rect 51548 1762 51604 3278
rect 51548 1710 51550 1762
rect 51602 1710 51604 1762
rect 51548 1698 51604 1710
rect 51772 3332 51828 3342
rect 51772 800 51828 3276
rect 52780 3332 52836 3342
rect 52780 3238 52836 3276
rect 53116 3332 53172 3342
rect 52444 1762 52500 1774
rect 52444 1710 52446 1762
rect 52498 1710 52500 1762
rect 52444 800 52500 1710
rect 53116 800 53172 3276
rect 53452 3330 53508 3342
rect 53452 3278 53454 3330
rect 53506 3278 53508 3330
rect 53452 1762 53508 3278
rect 54124 3332 54180 3342
rect 54124 3238 54180 3276
rect 54460 3332 54516 3342
rect 53452 1710 53454 1762
rect 53506 1710 53508 1762
rect 53452 1698 53508 1710
rect 53788 1762 53844 1774
rect 53788 1710 53790 1762
rect 53842 1710 53844 1762
rect 53788 800 53844 1710
rect 54460 800 54516 3276
rect 54796 3330 54852 3342
rect 54796 3278 54798 3330
rect 54850 3278 54852 3330
rect 54796 1762 54852 3278
rect 54796 1710 54798 1762
rect 54850 1710 54852 1762
rect 54796 1698 54852 1710
rect 55132 800 55188 4396
rect 55356 4386 55412 4396
rect 59164 4450 59444 4452
rect 59164 4398 59390 4450
rect 59442 4398 59444 4450
rect 59164 4396 59444 4398
rect 55468 3332 55524 3342
rect 55468 3238 55524 3276
rect 56476 3332 56532 3342
rect 55804 1762 55860 1774
rect 55804 1710 55806 1762
rect 55858 1710 55860 1762
rect 55804 800 55860 1710
rect 56476 800 56532 3276
rect 56700 3330 56756 3342
rect 56700 3278 56702 3330
rect 56754 3278 56756 3330
rect 56700 1762 56756 3278
rect 57372 3332 57428 3342
rect 57372 3238 57428 3276
rect 58044 3330 58100 3342
rect 58044 3278 58046 3330
rect 58098 3278 58100 3330
rect 57820 1874 57876 1886
rect 57820 1822 57822 1874
rect 57874 1822 57876 1874
rect 56700 1710 56702 1762
rect 56754 1710 56756 1762
rect 56700 1698 56756 1710
rect 57148 1762 57204 1774
rect 57148 1710 57150 1762
rect 57202 1710 57204 1762
rect 57148 800 57204 1710
rect 57820 800 57876 1822
rect 58044 1762 58100 3278
rect 58044 1710 58046 1762
rect 58098 1710 58100 1762
rect 58044 1698 58100 1710
rect 58492 3332 58548 3342
rect 58492 800 58548 3276
rect 58716 3330 58772 3342
rect 58716 3278 58718 3330
rect 58770 3278 58772 3330
rect 58716 1874 58772 3278
rect 58716 1822 58718 1874
rect 58770 1822 58772 1874
rect 58716 1810 58772 1822
rect 59164 800 59220 4396
rect 59388 4386 59444 4396
rect 63196 4450 63476 4452
rect 63196 4398 63422 4450
rect 63474 4398 63476 4450
rect 63196 4396 63476 4398
rect 59388 3332 59444 3342
rect 59388 3238 59444 3276
rect 59836 3332 59892 3342
rect 59836 800 59892 3276
rect 60620 3332 60676 3342
rect 60620 3238 60676 3276
rect 61292 3330 61348 3342
rect 61292 3278 61294 3330
rect 61346 3278 61348 3330
rect 61180 1874 61236 1886
rect 61180 1822 61182 1874
rect 61234 1822 61236 1874
rect 60508 1762 60564 1774
rect 60508 1710 60510 1762
rect 60562 1710 60564 1762
rect 60508 800 60564 1710
rect 61180 800 61236 1822
rect 61292 1762 61348 3278
rect 61292 1710 61294 1762
rect 61346 1710 61348 1762
rect 61292 1698 61348 1710
rect 61852 3332 61908 3342
rect 61852 800 61908 3276
rect 61964 3330 62020 3342
rect 61964 3278 61966 3330
rect 62018 3278 62020 3330
rect 61964 1874 62020 3278
rect 62636 3332 62692 3342
rect 62636 3238 62692 3276
rect 61964 1822 61966 1874
rect 62018 1822 62020 1874
rect 61964 1810 62020 1822
rect 62524 1762 62580 1774
rect 62524 1710 62526 1762
rect 62578 1710 62580 1762
rect 62524 800 62580 1710
rect 63196 800 63252 4396
rect 63420 4386 63476 4396
rect 70588 4450 70868 4452
rect 70588 4398 70814 4450
rect 70866 4398 70868 4450
rect 70588 4396 70868 4398
rect 65916 3948 66180 3958
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 65916 3882 66180 3892
rect 63308 3330 63364 3342
rect 63308 3278 63310 3330
rect 63362 3278 63364 3330
rect 63308 1762 63364 3278
rect 64540 3330 64596 3342
rect 64540 3278 64542 3330
rect 64594 3278 64596 3330
rect 63308 1710 63310 1762
rect 63362 1710 63364 1762
rect 63308 1698 63364 1710
rect 63868 1762 63924 1774
rect 63868 1710 63870 1762
rect 63922 1710 63924 1762
rect 63868 800 63924 1710
rect 64540 1762 64596 3278
rect 65212 3330 65268 3342
rect 65212 3278 65214 3330
rect 65266 3278 65268 3330
rect 64540 1710 64542 1762
rect 64594 1710 64596 1762
rect 64540 1698 64596 1710
rect 64652 1874 64708 1886
rect 64652 1822 64654 1874
rect 64706 1822 64708 1874
rect 64652 1540 64708 1822
rect 65212 1874 65268 3278
rect 65212 1822 65214 1874
rect 65266 1822 65268 1874
rect 65212 1810 65268 1822
rect 65324 3332 65380 3342
rect 65324 1540 65380 3276
rect 65884 3332 65940 3342
rect 65884 3238 65940 3276
rect 66556 3330 66612 3342
rect 66556 3278 66558 3330
rect 66610 3278 66612 3330
rect 64540 1484 64708 1540
rect 65212 1484 65380 1540
rect 65884 1874 65940 1886
rect 65884 1822 65886 1874
rect 65938 1822 65940 1874
rect 64540 800 64596 1484
rect 65212 800 65268 1484
rect 65884 800 65940 1822
rect 66556 1874 66612 3278
rect 66556 1822 66558 1874
rect 66610 1822 66612 1874
rect 66556 1810 66612 1822
rect 66668 3332 66724 3342
rect 66668 1652 66724 3276
rect 67228 3332 67284 3342
rect 67228 3238 67284 3276
rect 67900 3332 67956 3342
rect 66556 1596 66724 1652
rect 67228 1762 67284 1774
rect 67228 1710 67230 1762
rect 67282 1710 67284 1762
rect 66556 800 66612 1596
rect 67228 800 67284 1710
rect 67900 800 67956 3276
rect 68460 3330 68516 3342
rect 68460 3278 68462 3330
rect 68514 3278 68516 3330
rect 68460 1762 68516 3278
rect 69132 3332 69188 3342
rect 69132 3238 69188 3276
rect 69804 3330 69860 3342
rect 69804 3278 69806 3330
rect 69858 3278 69860 3330
rect 68460 1710 68462 1762
rect 68514 1710 68516 1762
rect 68460 1698 68516 1710
rect 68572 1764 68628 1774
rect 68572 800 68628 1708
rect 69244 1762 69300 1774
rect 69244 1710 69246 1762
rect 69298 1710 69300 1762
rect 69244 800 69300 1710
rect 69804 1764 69860 3278
rect 70476 3330 70532 3342
rect 70476 3278 70478 3330
rect 70530 3278 70532 3330
rect 69804 1698 69860 1708
rect 69916 1876 69972 1886
rect 69916 800 69972 1820
rect 70476 1762 70532 3278
rect 70476 1710 70478 1762
rect 70530 1710 70532 1762
rect 70476 1698 70532 1710
rect 70588 800 70644 4396
rect 70812 4386 70868 4396
rect 73164 4450 73444 4452
rect 73164 4398 73390 4450
rect 73442 4398 73444 4450
rect 73164 4396 73444 4398
rect 71148 3330 71204 3342
rect 71148 3278 71150 3330
rect 71202 3278 71204 3330
rect 71148 1876 71204 3278
rect 71148 1810 71204 1820
rect 71260 3332 71316 3342
rect 71260 800 71316 3276
rect 72380 3332 72436 3342
rect 72380 3238 72436 3276
rect 73052 3330 73108 3342
rect 73052 3278 73054 3330
rect 73106 3278 73108 3330
rect 71932 1764 71988 1774
rect 71932 800 71988 1708
rect 72604 1762 72660 1774
rect 72604 1710 72606 1762
rect 72658 1710 72660 1762
rect 72604 800 72660 1710
rect 73052 1764 73108 3278
rect 73052 1698 73108 1708
rect 73164 1540 73220 4396
rect 73388 4386 73444 4396
rect 73500 4452 73556 4462
rect 73052 1484 73220 1540
rect 73276 3332 73332 3342
rect 73052 800 73108 1484
rect 73276 800 73332 3276
rect 73500 800 73556 4396
rect 74060 4452 74116 4462
rect 74060 4358 74116 4396
rect 73724 3330 73780 3342
rect 73724 3278 73726 3330
rect 73778 3278 73780 3330
rect 73724 1762 73780 3278
rect 74396 3332 74452 3342
rect 74396 3238 74452 3276
rect 73724 1710 73726 1762
rect 73778 1710 73780 1762
rect 73724 1698 73780 1710
rect 6272 0 6384 800
rect 6496 0 6608 800
rect 6720 0 6832 800
rect 6944 0 7056 800
rect 7168 0 7280 800
rect 7392 0 7504 800
rect 7616 0 7728 800
rect 7840 0 7952 800
rect 8064 0 8176 800
rect 8288 0 8400 800
rect 8512 0 8624 800
rect 8736 0 8848 800
rect 8960 0 9072 800
rect 9184 0 9296 800
rect 9408 0 9520 800
rect 9632 0 9744 800
rect 9856 0 9968 800
rect 10080 0 10192 800
rect 10304 0 10416 800
rect 10528 0 10640 800
rect 10752 0 10864 800
rect 10976 0 11088 800
rect 11200 0 11312 800
rect 11424 0 11536 800
rect 11648 0 11760 800
rect 11872 0 11984 800
rect 12096 0 12208 800
rect 12320 0 12432 800
rect 12544 0 12656 800
rect 12768 0 12880 800
rect 12992 0 13104 800
rect 13216 0 13328 800
rect 13440 0 13552 800
rect 13664 0 13776 800
rect 13888 0 14000 800
rect 14112 0 14224 800
rect 14336 0 14448 800
rect 14560 0 14672 800
rect 14784 0 14896 800
rect 15008 0 15120 800
rect 15232 0 15344 800
rect 15456 0 15568 800
rect 15680 0 15792 800
rect 15904 0 16016 800
rect 16128 0 16240 800
rect 16352 0 16464 800
rect 16576 0 16688 800
rect 16800 0 16912 800
rect 17024 0 17136 800
rect 17248 0 17360 800
rect 17472 0 17584 800
rect 17696 0 17808 800
rect 17920 0 18032 800
rect 18144 0 18256 800
rect 18368 0 18480 800
rect 18592 0 18704 800
rect 18816 0 18928 800
rect 19040 0 19152 800
rect 19264 0 19376 800
rect 19488 0 19600 800
rect 19712 0 19824 800
rect 19936 0 20048 800
rect 20160 0 20272 800
rect 20384 0 20496 800
rect 20608 0 20720 800
rect 20832 0 20944 800
rect 21056 0 21168 800
rect 21280 0 21392 800
rect 21504 0 21616 800
rect 21728 0 21840 800
rect 21952 0 22064 800
rect 22176 0 22288 800
rect 22400 0 22512 800
rect 22624 0 22736 800
rect 22848 0 22960 800
rect 23072 0 23184 800
rect 23296 0 23408 800
rect 23520 0 23632 800
rect 23744 0 23856 800
rect 23968 0 24080 800
rect 24192 0 24304 800
rect 24416 0 24528 800
rect 24640 0 24752 800
rect 24864 0 24976 800
rect 25088 0 25200 800
rect 25312 0 25424 800
rect 25536 0 25648 800
rect 25760 0 25872 800
rect 25984 0 26096 800
rect 26208 0 26320 800
rect 26432 0 26544 800
rect 26656 0 26768 800
rect 26880 0 26992 800
rect 27104 0 27216 800
rect 27328 0 27440 800
rect 27552 0 27664 800
rect 27776 0 27888 800
rect 28000 0 28112 800
rect 28224 0 28336 800
rect 28448 0 28560 800
rect 28672 0 28784 800
rect 28896 0 29008 800
rect 29120 0 29232 800
rect 29344 0 29456 800
rect 29568 0 29680 800
rect 29792 0 29904 800
rect 30016 0 30128 800
rect 30240 0 30352 800
rect 30464 0 30576 800
rect 30688 0 30800 800
rect 30912 0 31024 800
rect 31136 0 31248 800
rect 31360 0 31472 800
rect 31584 0 31696 800
rect 31808 0 31920 800
rect 32032 0 32144 800
rect 32256 0 32368 800
rect 32480 0 32592 800
rect 32704 0 32816 800
rect 32928 0 33040 800
rect 33152 0 33264 800
rect 33376 0 33488 800
rect 33600 0 33712 800
rect 33824 0 33936 800
rect 34048 0 34160 800
rect 34272 0 34384 800
rect 34496 0 34608 800
rect 34720 0 34832 800
rect 34944 0 35056 800
rect 35168 0 35280 800
rect 35392 0 35504 800
rect 35616 0 35728 800
rect 35840 0 35952 800
rect 36064 0 36176 800
rect 36288 0 36400 800
rect 36512 0 36624 800
rect 36736 0 36848 800
rect 36960 0 37072 800
rect 37184 0 37296 800
rect 37408 0 37520 800
rect 37632 0 37744 800
rect 37856 0 37968 800
rect 38080 0 38192 800
rect 38304 0 38416 800
rect 38528 0 38640 800
rect 38752 0 38864 800
rect 38976 0 39088 800
rect 39200 0 39312 800
rect 39424 0 39536 800
rect 39648 0 39760 800
rect 39872 0 39984 800
rect 40096 0 40208 800
rect 40320 0 40432 800
rect 40544 0 40656 800
rect 40768 0 40880 800
rect 40992 0 41104 800
rect 41216 0 41328 800
rect 41440 0 41552 800
rect 41664 0 41776 800
rect 41888 0 42000 800
rect 42112 0 42224 800
rect 42336 0 42448 800
rect 42560 0 42672 800
rect 42784 0 42896 800
rect 43008 0 43120 800
rect 43232 0 43344 800
rect 43456 0 43568 800
rect 43680 0 43792 800
rect 43904 0 44016 800
rect 44128 0 44240 800
rect 44352 0 44464 800
rect 44576 0 44688 800
rect 44800 0 44912 800
rect 45024 0 45136 800
rect 45248 0 45360 800
rect 45472 0 45584 800
rect 45696 0 45808 800
rect 45920 0 46032 800
rect 46144 0 46256 800
rect 46368 0 46480 800
rect 46592 0 46704 800
rect 46816 0 46928 800
rect 47040 0 47152 800
rect 47264 0 47376 800
rect 47488 0 47600 800
rect 47712 0 47824 800
rect 47936 0 48048 800
rect 48160 0 48272 800
rect 48384 0 48496 800
rect 48608 0 48720 800
rect 48832 0 48944 800
rect 49056 0 49168 800
rect 49280 0 49392 800
rect 49504 0 49616 800
rect 49728 0 49840 800
rect 49952 0 50064 800
rect 50176 0 50288 800
rect 50400 0 50512 800
rect 50624 0 50736 800
rect 50848 0 50960 800
rect 51072 0 51184 800
rect 51296 0 51408 800
rect 51520 0 51632 800
rect 51744 0 51856 800
rect 51968 0 52080 800
rect 52192 0 52304 800
rect 52416 0 52528 800
rect 52640 0 52752 800
rect 52864 0 52976 800
rect 53088 0 53200 800
rect 53312 0 53424 800
rect 53536 0 53648 800
rect 53760 0 53872 800
rect 53984 0 54096 800
rect 54208 0 54320 800
rect 54432 0 54544 800
rect 54656 0 54768 800
rect 54880 0 54992 800
rect 55104 0 55216 800
rect 55328 0 55440 800
rect 55552 0 55664 800
rect 55776 0 55888 800
rect 56000 0 56112 800
rect 56224 0 56336 800
rect 56448 0 56560 800
rect 56672 0 56784 800
rect 56896 0 57008 800
rect 57120 0 57232 800
rect 57344 0 57456 800
rect 57568 0 57680 800
rect 57792 0 57904 800
rect 58016 0 58128 800
rect 58240 0 58352 800
rect 58464 0 58576 800
rect 58688 0 58800 800
rect 58912 0 59024 800
rect 59136 0 59248 800
rect 59360 0 59472 800
rect 59584 0 59696 800
rect 59808 0 59920 800
rect 60032 0 60144 800
rect 60256 0 60368 800
rect 60480 0 60592 800
rect 60704 0 60816 800
rect 60928 0 61040 800
rect 61152 0 61264 800
rect 61376 0 61488 800
rect 61600 0 61712 800
rect 61824 0 61936 800
rect 62048 0 62160 800
rect 62272 0 62384 800
rect 62496 0 62608 800
rect 62720 0 62832 800
rect 62944 0 63056 800
rect 63168 0 63280 800
rect 63392 0 63504 800
rect 63616 0 63728 800
rect 63840 0 63952 800
rect 64064 0 64176 800
rect 64288 0 64400 800
rect 64512 0 64624 800
rect 64736 0 64848 800
rect 64960 0 65072 800
rect 65184 0 65296 800
rect 65408 0 65520 800
rect 65632 0 65744 800
rect 65856 0 65968 800
rect 66080 0 66192 800
rect 66304 0 66416 800
rect 66528 0 66640 800
rect 66752 0 66864 800
rect 66976 0 67088 800
rect 67200 0 67312 800
rect 67424 0 67536 800
rect 67648 0 67760 800
rect 67872 0 67984 800
rect 68096 0 68208 800
rect 68320 0 68432 800
rect 68544 0 68656 800
rect 68768 0 68880 800
rect 68992 0 69104 800
rect 69216 0 69328 800
rect 69440 0 69552 800
rect 69664 0 69776 800
rect 69888 0 70000 800
rect 70112 0 70224 800
rect 70336 0 70448 800
rect 70560 0 70672 800
rect 70784 0 70896 800
rect 71008 0 71120 800
rect 71232 0 71344 800
rect 71456 0 71568 800
rect 71680 0 71792 800
rect 71904 0 72016 800
rect 72128 0 72240 800
rect 72352 0 72464 800
rect 72576 0 72688 800
rect 72800 0 72912 800
rect 73024 0 73136 800
rect 73248 0 73360 800
rect 73472 0 73584 800
<< via2 >>
rect 2940 76636 2996 76692
rect 3836 76690 3892 76692
rect 3836 76638 3838 76690
rect 3838 76638 3890 76690
rect 3890 76638 3892 76690
rect 3836 76636 3892 76638
rect 3612 76524 3668 76580
rect 4476 76074 4532 76076
rect 4476 76022 4478 76074
rect 4478 76022 4530 76074
rect 4530 76022 4532 76074
rect 4476 76020 4532 76022
rect 4580 76074 4636 76076
rect 4580 76022 4582 76074
rect 4582 76022 4634 76074
rect 4634 76022 4636 76074
rect 4580 76020 4636 76022
rect 4684 76074 4740 76076
rect 4684 76022 4686 76074
rect 4686 76022 4738 76074
rect 4738 76022 4740 76074
rect 4684 76020 4740 76022
rect 3388 75852 3444 75908
rect 6860 76636 6916 76692
rect 5852 76578 5908 76580
rect 5852 76526 5854 76578
rect 5854 76526 5906 76578
rect 5906 76526 5908 76578
rect 5852 76524 5908 76526
rect 7980 76636 8036 76692
rect 4476 74506 4532 74508
rect 4476 74454 4478 74506
rect 4478 74454 4530 74506
rect 4530 74454 4532 74506
rect 4476 74452 4532 74454
rect 4580 74506 4636 74508
rect 4580 74454 4582 74506
rect 4582 74454 4634 74506
rect 4634 74454 4636 74506
rect 4580 74452 4636 74454
rect 4684 74506 4740 74508
rect 4684 74454 4686 74506
rect 4686 74454 4738 74506
rect 4738 74454 4740 74506
rect 4684 74452 4740 74454
rect 4476 72938 4532 72940
rect 4476 72886 4478 72938
rect 4478 72886 4530 72938
rect 4530 72886 4532 72938
rect 4476 72884 4532 72886
rect 4580 72938 4636 72940
rect 4580 72886 4582 72938
rect 4582 72886 4634 72938
rect 4634 72886 4636 72938
rect 4580 72884 4636 72886
rect 4684 72938 4740 72940
rect 4684 72886 4686 72938
rect 4686 72886 4738 72938
rect 4738 72886 4740 72938
rect 4684 72884 4740 72886
rect 14924 76466 14980 76468
rect 14924 76414 14926 76466
rect 14926 76414 14978 76466
rect 14978 76414 14980 76466
rect 14924 76412 14980 76414
rect 13020 75516 13076 75572
rect 13692 75570 13748 75572
rect 13692 75518 13694 75570
rect 13694 75518 13746 75570
rect 13746 75518 13748 75570
rect 13692 75516 13748 75518
rect 15820 76412 15876 76468
rect 16716 75628 16772 75684
rect 18844 76466 18900 76468
rect 18844 76414 18846 76466
rect 18846 76414 18898 76466
rect 18898 76414 18900 76466
rect 18844 76412 18900 76414
rect 17836 75682 17892 75684
rect 17836 75630 17838 75682
rect 17838 75630 17890 75682
rect 17890 75630 17892 75682
rect 17836 75628 17892 75630
rect 19836 76858 19892 76860
rect 19836 76806 19838 76858
rect 19838 76806 19890 76858
rect 19890 76806 19892 76858
rect 19836 76804 19892 76806
rect 19940 76858 19996 76860
rect 19940 76806 19942 76858
rect 19942 76806 19994 76858
rect 19994 76806 19996 76858
rect 19940 76804 19996 76806
rect 20044 76858 20100 76860
rect 20044 76806 20046 76858
rect 20046 76806 20098 76858
rect 20098 76806 20100 76858
rect 20044 76804 20100 76806
rect 19852 76412 19908 76468
rect 19852 76188 19908 76244
rect 20860 75964 20916 76020
rect 21756 75852 21812 75908
rect 21084 75516 21140 75572
rect 21644 75570 21700 75572
rect 21644 75518 21646 75570
rect 21646 75518 21698 75570
rect 21698 75518 21700 75570
rect 21644 75516 21700 75518
rect 15820 75404 15876 75460
rect 21420 75404 21476 75460
rect 19836 75290 19892 75292
rect 19836 75238 19838 75290
rect 19838 75238 19890 75290
rect 19890 75238 19892 75290
rect 19836 75236 19892 75238
rect 19940 75290 19996 75292
rect 19940 75238 19942 75290
rect 19942 75238 19994 75290
rect 19994 75238 19996 75290
rect 19940 75236 19996 75238
rect 20044 75290 20100 75292
rect 20044 75238 20046 75290
rect 20046 75238 20098 75290
rect 20098 75238 20100 75290
rect 20044 75236 20100 75238
rect 19836 73722 19892 73724
rect 19836 73670 19838 73722
rect 19838 73670 19890 73722
rect 19890 73670 19892 73722
rect 19836 73668 19892 73670
rect 19940 73722 19996 73724
rect 19940 73670 19942 73722
rect 19942 73670 19994 73722
rect 19994 73670 19996 73722
rect 19940 73668 19996 73670
rect 20044 73722 20100 73724
rect 20044 73670 20046 73722
rect 20046 73670 20098 73722
rect 20098 73670 20100 73722
rect 20044 73668 20100 73670
rect 12908 72492 12964 72548
rect 22764 75852 22820 75908
rect 23996 75852 24052 75908
rect 24780 75794 24836 75796
rect 24780 75742 24782 75794
rect 24782 75742 24834 75794
rect 24834 75742 24836 75794
rect 24780 75740 24836 75742
rect 28476 75740 28532 75796
rect 27916 75570 27972 75572
rect 27916 75518 27918 75570
rect 27918 75518 27970 75570
rect 27970 75518 27972 75570
rect 27916 75516 27972 75518
rect 28140 75404 28196 75460
rect 26572 74396 26628 74452
rect 21756 74284 21812 74340
rect 29148 75740 29204 75796
rect 29932 75516 29988 75572
rect 30044 75628 30100 75684
rect 28588 74172 28644 74228
rect 28812 74284 28868 74340
rect 30156 75404 30212 75460
rect 30492 75404 30548 75460
rect 30268 75122 30324 75124
rect 30268 75070 30270 75122
rect 30270 75070 30322 75122
rect 30322 75070 30324 75122
rect 30268 75068 30324 75070
rect 29372 74284 29428 74340
rect 29708 74226 29764 74228
rect 29708 74174 29710 74226
rect 29710 74174 29762 74226
rect 29762 74174 29764 74226
rect 29708 74172 29764 74174
rect 28812 73948 28868 74004
rect 29484 73948 29540 74004
rect 30156 74002 30212 74004
rect 30156 73950 30158 74002
rect 30158 73950 30210 74002
rect 30210 73950 30212 74002
rect 30156 73948 30212 73950
rect 30940 75682 30996 75684
rect 30940 75630 30942 75682
rect 30942 75630 30994 75682
rect 30994 75630 30996 75682
rect 30940 75628 30996 75630
rect 30716 75292 30772 75348
rect 30940 75180 30996 75236
rect 31500 75404 31556 75460
rect 31164 75180 31220 75236
rect 30716 74898 30772 74900
rect 30716 74846 30718 74898
rect 30718 74846 30770 74898
rect 30770 74846 30772 74898
rect 30716 74844 30772 74846
rect 31500 75068 31556 75124
rect 31164 74172 31220 74228
rect 31052 74002 31108 74004
rect 31052 73950 31054 74002
rect 31054 73950 31106 74002
rect 31106 73950 31108 74002
rect 31052 73948 31108 73950
rect 31388 73890 31444 73892
rect 31388 73838 31390 73890
rect 31390 73838 31442 73890
rect 31442 73838 31444 73890
rect 31388 73836 31444 73838
rect 28476 73388 28532 73444
rect 30940 73388 30996 73444
rect 30380 72716 30436 72772
rect 31276 73442 31332 73444
rect 31276 73390 31278 73442
rect 31278 73390 31330 73442
rect 31330 73390 31332 73442
rect 31276 73388 31332 73390
rect 31836 75740 31892 75796
rect 32060 75068 32116 75124
rect 32060 74844 32116 74900
rect 31948 74396 32004 74452
rect 32732 75794 32788 75796
rect 32732 75742 32734 75794
rect 32734 75742 32786 75794
rect 32786 75742 32788 75794
rect 32732 75740 32788 75742
rect 34412 77644 34468 77700
rect 34300 76188 34356 76244
rect 34188 75964 34244 76020
rect 33180 75516 33236 75572
rect 32844 75404 32900 75460
rect 32620 74786 32676 74788
rect 32620 74734 32622 74786
rect 32622 74734 32674 74786
rect 32674 74734 32676 74786
rect 32620 74732 32676 74734
rect 32620 74396 32676 74452
rect 32172 74226 32228 74228
rect 32172 74174 32174 74226
rect 32174 74174 32226 74226
rect 32226 74174 32228 74226
rect 32172 74172 32228 74174
rect 31612 73500 31668 73556
rect 21420 72380 21476 72436
rect 32060 73554 32116 73556
rect 32060 73502 32062 73554
rect 32062 73502 32114 73554
rect 32114 73502 32116 73554
rect 32060 73500 32116 73502
rect 33068 75068 33124 75124
rect 33740 75010 33796 75012
rect 33740 74958 33742 75010
rect 33742 74958 33794 75010
rect 33794 74958 33796 75010
rect 33740 74956 33796 74958
rect 32620 73500 32676 73556
rect 32956 73612 33012 73668
rect 34412 75068 34468 75124
rect 35644 77532 35700 77588
rect 34076 74732 34132 74788
rect 34188 74338 34244 74340
rect 34188 74286 34190 74338
rect 34190 74286 34242 74338
rect 34242 74286 34244 74338
rect 34188 74284 34244 74286
rect 33852 74172 33908 74228
rect 34300 74172 34356 74228
rect 33292 73836 33348 73892
rect 33740 73612 33796 73668
rect 33628 73554 33684 73556
rect 33628 73502 33630 73554
rect 33630 73502 33682 73554
rect 33682 73502 33684 73554
rect 33628 73500 33684 73502
rect 33404 73388 33460 73444
rect 19836 72154 19892 72156
rect 19836 72102 19838 72154
rect 19838 72102 19890 72154
rect 19890 72102 19892 72154
rect 19836 72100 19892 72102
rect 19940 72154 19996 72156
rect 19940 72102 19942 72154
rect 19942 72102 19994 72154
rect 19994 72102 19996 72154
rect 19940 72100 19996 72102
rect 20044 72154 20100 72156
rect 20044 72102 20046 72154
rect 20046 72102 20098 72154
rect 20098 72102 20100 72154
rect 20044 72100 20100 72102
rect 4476 71370 4532 71372
rect 4476 71318 4478 71370
rect 4478 71318 4530 71370
rect 4530 71318 4532 71370
rect 4476 71316 4532 71318
rect 4580 71370 4636 71372
rect 4580 71318 4582 71370
rect 4582 71318 4634 71370
rect 4634 71318 4636 71370
rect 4580 71316 4636 71318
rect 4684 71370 4740 71372
rect 4684 71318 4686 71370
rect 4686 71318 4738 71370
rect 4738 71318 4740 71370
rect 4684 71316 4740 71318
rect 19836 70586 19892 70588
rect 19836 70534 19838 70586
rect 19838 70534 19890 70586
rect 19890 70534 19892 70586
rect 19836 70532 19892 70534
rect 19940 70586 19996 70588
rect 19940 70534 19942 70586
rect 19942 70534 19994 70586
rect 19994 70534 19996 70586
rect 19940 70532 19996 70534
rect 20044 70586 20100 70588
rect 20044 70534 20046 70586
rect 20046 70534 20098 70586
rect 20098 70534 20100 70586
rect 20044 70532 20100 70534
rect 34524 74898 34580 74900
rect 34524 74846 34526 74898
rect 34526 74846 34578 74898
rect 34578 74846 34580 74898
rect 34524 74844 34580 74846
rect 34524 74226 34580 74228
rect 34524 74174 34526 74226
rect 34526 74174 34578 74226
rect 34578 74174 34580 74226
rect 34524 74172 34580 74174
rect 34636 73948 34692 74004
rect 34748 74114 34804 74116
rect 34748 74062 34750 74114
rect 34750 74062 34802 74114
rect 34802 74062 34804 74114
rect 34748 74060 34804 74062
rect 34412 73612 34468 73668
rect 34524 73442 34580 73444
rect 34524 73390 34526 73442
rect 34526 73390 34578 73442
rect 34578 73390 34580 73442
rect 34524 73388 34580 73390
rect 35196 76074 35252 76076
rect 35196 76022 35198 76074
rect 35198 76022 35250 76074
rect 35250 76022 35252 76074
rect 35196 76020 35252 76022
rect 35300 76074 35356 76076
rect 35300 76022 35302 76074
rect 35302 76022 35354 76074
rect 35354 76022 35356 76074
rect 35300 76020 35356 76022
rect 35404 76074 35460 76076
rect 35404 76022 35406 76074
rect 35406 76022 35458 76074
rect 35458 76022 35460 76074
rect 35404 76020 35460 76022
rect 36092 75964 36148 76020
rect 36204 75852 36260 75908
rect 35756 75068 35812 75124
rect 35196 74506 35252 74508
rect 35196 74454 35198 74506
rect 35198 74454 35250 74506
rect 35250 74454 35252 74506
rect 35196 74452 35252 74454
rect 35300 74506 35356 74508
rect 35300 74454 35302 74506
rect 35302 74454 35354 74506
rect 35354 74454 35356 74506
rect 35300 74452 35356 74454
rect 35404 74506 35460 74508
rect 35404 74454 35406 74506
rect 35406 74454 35458 74506
rect 35458 74454 35460 74506
rect 35404 74452 35460 74454
rect 35644 74844 35700 74900
rect 35644 74396 35700 74452
rect 35308 74172 35364 74228
rect 35420 74002 35476 74004
rect 35420 73950 35422 74002
rect 35422 73950 35474 74002
rect 35474 73950 35476 74002
rect 35420 73948 35476 73950
rect 36092 74844 36148 74900
rect 35980 74114 36036 74116
rect 35980 74062 35982 74114
rect 35982 74062 36034 74114
rect 36034 74062 36036 74114
rect 35980 74060 36036 74062
rect 35196 72938 35252 72940
rect 35196 72886 35198 72938
rect 35198 72886 35250 72938
rect 35250 72886 35252 72938
rect 35196 72884 35252 72886
rect 35300 72938 35356 72940
rect 35300 72886 35302 72938
rect 35302 72886 35354 72938
rect 35354 72886 35356 72938
rect 35300 72884 35356 72886
rect 35404 72938 35460 72940
rect 35404 72886 35406 72938
rect 35406 72886 35458 72938
rect 35458 72886 35460 72938
rect 35404 72884 35460 72886
rect 35084 72546 35140 72548
rect 35084 72494 35086 72546
rect 35086 72494 35138 72546
rect 35138 72494 35140 72546
rect 35084 72492 35140 72494
rect 34412 72434 34468 72436
rect 34412 72382 34414 72434
rect 34414 72382 34466 72434
rect 34466 72382 34468 72434
rect 34412 72380 34468 72382
rect 35196 72434 35252 72436
rect 35196 72382 35198 72434
rect 35198 72382 35250 72434
rect 35250 72382 35252 72434
rect 35196 72380 35252 72382
rect 36428 74732 36484 74788
rect 36204 72604 36260 72660
rect 36204 72380 36260 72436
rect 34748 71874 34804 71876
rect 34748 71822 34750 71874
rect 34750 71822 34802 71874
rect 34802 71822 34804 71874
rect 34748 71820 34804 71822
rect 35196 71370 35252 71372
rect 35196 71318 35198 71370
rect 35198 71318 35250 71370
rect 35250 71318 35252 71370
rect 35196 71316 35252 71318
rect 35300 71370 35356 71372
rect 35300 71318 35302 71370
rect 35302 71318 35354 71370
rect 35354 71318 35356 71370
rect 35300 71316 35356 71318
rect 35404 71370 35460 71372
rect 35404 71318 35406 71370
rect 35406 71318 35458 71370
rect 35458 71318 35460 71370
rect 35404 71316 35460 71318
rect 34300 71036 34356 71092
rect 35308 71090 35364 71092
rect 35308 71038 35310 71090
rect 35310 71038 35362 71090
rect 35362 71038 35364 71090
rect 35308 71036 35364 71038
rect 31948 70476 32004 70532
rect 36540 74284 36596 74340
rect 37212 76412 37268 76468
rect 37100 76300 37156 76356
rect 37884 76354 37940 76356
rect 37884 76302 37886 76354
rect 37886 76302 37938 76354
rect 37938 76302 37940 76354
rect 37884 76300 37940 76302
rect 37212 76242 37268 76244
rect 37212 76190 37214 76242
rect 37214 76190 37266 76242
rect 37266 76190 37268 76242
rect 37212 76188 37268 76190
rect 38556 76524 38612 76580
rect 36988 74844 37044 74900
rect 36764 74508 36820 74564
rect 36652 73500 36708 73556
rect 36988 74508 37044 74564
rect 36876 73836 36932 73892
rect 36540 72716 36596 72772
rect 36540 72434 36596 72436
rect 36540 72382 36542 72434
rect 36542 72382 36594 72434
rect 36594 72382 36596 72434
rect 36540 72380 36596 72382
rect 36428 72268 36484 72324
rect 36876 72268 36932 72324
rect 36428 72044 36484 72100
rect 36876 71260 36932 71316
rect 36428 71090 36484 71092
rect 36428 71038 36430 71090
rect 36430 71038 36482 71090
rect 36482 71038 36484 71090
rect 36428 71036 36484 71038
rect 36316 70364 36372 70420
rect 37100 70418 37156 70420
rect 37100 70366 37102 70418
rect 37102 70366 37154 70418
rect 37154 70366 37156 70418
rect 37100 70364 37156 70366
rect 37660 75458 37716 75460
rect 37660 75406 37662 75458
rect 37662 75406 37714 75458
rect 37714 75406 37716 75458
rect 37660 75404 37716 75406
rect 37548 74114 37604 74116
rect 37548 74062 37550 74114
rect 37550 74062 37602 74114
rect 37602 74062 37604 74114
rect 37548 74060 37604 74062
rect 37884 74844 37940 74900
rect 37772 74060 37828 74116
rect 37548 73276 37604 73332
rect 37996 74508 38052 74564
rect 38108 74060 38164 74116
rect 37996 73724 38052 73780
rect 38444 74898 38500 74900
rect 38444 74846 38446 74898
rect 38446 74846 38498 74898
rect 38498 74846 38500 74898
rect 38444 74844 38500 74846
rect 38892 76578 38948 76580
rect 38892 76526 38894 76578
rect 38894 76526 38946 76578
rect 38946 76526 38948 76578
rect 38892 76524 38948 76526
rect 39564 76300 39620 76356
rect 39452 76188 39508 76244
rect 38780 75010 38836 75012
rect 38780 74958 38782 75010
rect 38782 74958 38834 75010
rect 38834 74958 38836 75010
rect 38780 74956 38836 74958
rect 38892 74844 38948 74900
rect 39452 75740 39508 75796
rect 39004 74002 39060 74004
rect 39004 73950 39006 74002
rect 39006 73950 39058 74002
rect 39058 73950 39060 74002
rect 39004 73948 39060 73950
rect 38220 73612 38276 73668
rect 38220 73330 38276 73332
rect 38220 73278 38222 73330
rect 38222 73278 38274 73330
rect 38274 73278 38276 73330
rect 38220 73276 38276 73278
rect 37436 72434 37492 72436
rect 37436 72382 37438 72434
rect 37438 72382 37490 72434
rect 37490 72382 37492 72434
rect 37436 72380 37492 72382
rect 37660 72156 37716 72212
rect 37324 71932 37380 71988
rect 37548 72044 37604 72100
rect 37436 70306 37492 70308
rect 37436 70254 37438 70306
rect 37438 70254 37490 70306
rect 37490 70254 37492 70306
rect 37436 70252 37492 70254
rect 37212 70140 37268 70196
rect 37772 72044 37828 72100
rect 37884 72380 37940 72436
rect 37996 72156 38052 72212
rect 38332 71932 38388 71988
rect 38108 70866 38164 70868
rect 38108 70814 38110 70866
rect 38110 70814 38162 70866
rect 38162 70814 38164 70866
rect 38108 70812 38164 70814
rect 38668 73612 38724 73668
rect 38668 73330 38724 73332
rect 38668 73278 38670 73330
rect 38670 73278 38722 73330
rect 38722 73278 38724 73330
rect 38668 73276 38724 73278
rect 38556 72156 38612 72212
rect 39788 75628 39844 75684
rect 39676 75292 39732 75348
rect 40572 76524 40628 76580
rect 41132 76524 41188 76580
rect 40124 76412 40180 76468
rect 41020 76354 41076 76356
rect 41020 76302 41022 76354
rect 41022 76302 41074 76354
rect 41074 76302 41076 76354
rect 41020 76300 41076 76302
rect 40348 76188 40404 76244
rect 40012 75740 40068 75796
rect 40684 75682 40740 75684
rect 40684 75630 40686 75682
rect 40686 75630 40738 75682
rect 40738 75630 40740 75682
rect 40684 75628 40740 75630
rect 40796 75516 40852 75572
rect 40124 75180 40180 75236
rect 40236 75458 40292 75460
rect 40236 75406 40238 75458
rect 40238 75406 40290 75458
rect 40290 75406 40292 75458
rect 40236 75404 40292 75406
rect 39900 75068 39956 75124
rect 39676 74844 39732 74900
rect 40124 74226 40180 74228
rect 40124 74174 40126 74226
rect 40126 74174 40178 74226
rect 40178 74174 40180 74226
rect 40124 74172 40180 74174
rect 40460 74060 40516 74116
rect 38892 72434 38948 72436
rect 38892 72382 38894 72434
rect 38894 72382 38946 72434
rect 38946 72382 38948 72434
rect 38892 72380 38948 72382
rect 38780 72156 38836 72212
rect 38780 71148 38836 71204
rect 38556 70924 38612 70980
rect 38780 70812 38836 70868
rect 39116 72716 39172 72772
rect 40236 73724 40292 73780
rect 40572 74956 40628 75012
rect 40796 74956 40852 75012
rect 40572 73948 40628 74004
rect 40684 74284 40740 74340
rect 40572 73554 40628 73556
rect 40572 73502 40574 73554
rect 40574 73502 40626 73554
rect 40626 73502 40628 73554
rect 40572 73500 40628 73502
rect 40796 74114 40852 74116
rect 40796 74062 40798 74114
rect 40798 74062 40850 74114
rect 40850 74062 40852 74114
rect 40796 74060 40852 74062
rect 40460 73276 40516 73332
rect 40236 72716 40292 72772
rect 40124 71596 40180 71652
rect 39676 71202 39732 71204
rect 39676 71150 39678 71202
rect 39678 71150 39730 71202
rect 39730 71150 39732 71202
rect 39676 71148 39732 71150
rect 39676 70978 39732 70980
rect 39676 70926 39678 70978
rect 39678 70926 39730 70978
rect 39730 70926 39732 70978
rect 39676 70924 39732 70926
rect 40236 71036 40292 71092
rect 40012 70812 40068 70868
rect 40460 70812 40516 70868
rect 40348 70306 40404 70308
rect 40348 70254 40350 70306
rect 40350 70254 40402 70306
rect 40402 70254 40404 70306
rect 40348 70252 40404 70254
rect 40236 70194 40292 70196
rect 40236 70142 40238 70194
rect 40238 70142 40290 70194
rect 40290 70142 40292 70194
rect 40236 70140 40292 70142
rect 4476 69802 4532 69804
rect 4476 69750 4478 69802
rect 4478 69750 4530 69802
rect 4530 69750 4532 69802
rect 4476 69748 4532 69750
rect 4580 69802 4636 69804
rect 4580 69750 4582 69802
rect 4582 69750 4634 69802
rect 4634 69750 4636 69802
rect 4580 69748 4636 69750
rect 4684 69802 4740 69804
rect 4684 69750 4686 69802
rect 4686 69750 4738 69802
rect 4738 69750 4740 69802
rect 4684 69748 4740 69750
rect 35196 69802 35252 69804
rect 35196 69750 35198 69802
rect 35198 69750 35250 69802
rect 35250 69750 35252 69802
rect 35196 69748 35252 69750
rect 35300 69802 35356 69804
rect 35300 69750 35302 69802
rect 35302 69750 35354 69802
rect 35354 69750 35356 69802
rect 35300 69748 35356 69750
rect 35404 69802 35460 69804
rect 35404 69750 35406 69802
rect 35406 69750 35458 69802
rect 35458 69750 35460 69802
rect 35404 69748 35460 69750
rect 40796 70306 40852 70308
rect 40796 70254 40798 70306
rect 40798 70254 40850 70306
rect 40850 70254 40852 70306
rect 40796 70252 40852 70254
rect 41244 72156 41300 72212
rect 41244 71708 41300 71764
rect 41020 71090 41076 71092
rect 41020 71038 41022 71090
rect 41022 71038 41074 71090
rect 41074 71038 41076 71090
rect 41020 71036 41076 71038
rect 41692 76412 41748 76468
rect 41468 76188 41524 76244
rect 41692 76188 41748 76244
rect 41804 75570 41860 75572
rect 41804 75518 41806 75570
rect 41806 75518 41858 75570
rect 41858 75518 41860 75570
rect 41804 75516 41860 75518
rect 41692 74844 41748 74900
rect 42028 76578 42084 76580
rect 42028 76526 42030 76578
rect 42030 76526 42082 76578
rect 42082 76526 42084 76578
rect 42028 76524 42084 76526
rect 42588 76524 42644 76580
rect 43372 76690 43428 76692
rect 43372 76638 43374 76690
rect 43374 76638 43426 76690
rect 43426 76638 43428 76690
rect 43372 76636 43428 76638
rect 43036 76466 43092 76468
rect 43036 76414 43038 76466
rect 43038 76414 43090 76466
rect 43090 76414 43092 76466
rect 43036 76412 43092 76414
rect 42476 76076 42532 76132
rect 42252 75516 42308 75572
rect 41580 74060 41636 74116
rect 41468 73554 41524 73556
rect 41468 73502 41470 73554
rect 41470 73502 41522 73554
rect 41522 73502 41524 73554
rect 41468 73500 41524 73502
rect 42140 74396 42196 74452
rect 41804 73948 41860 74004
rect 42252 74284 42308 74340
rect 41916 73724 41972 73780
rect 41804 72940 41860 72996
rect 41580 72546 41636 72548
rect 41580 72494 41582 72546
rect 41582 72494 41634 72546
rect 41634 72494 41636 72546
rect 41580 72492 41636 72494
rect 41468 72322 41524 72324
rect 41468 72270 41470 72322
rect 41470 72270 41522 72322
rect 41522 72270 41524 72322
rect 41468 72268 41524 72270
rect 41692 72268 41748 72324
rect 41804 72380 41860 72436
rect 41916 72156 41972 72212
rect 41916 71596 41972 71652
rect 42364 74844 42420 74900
rect 42364 73388 42420 73444
rect 43036 75682 43092 75684
rect 43036 75630 43038 75682
rect 43038 75630 43090 75682
rect 43090 75630 43092 75682
rect 43036 75628 43092 75630
rect 42812 75570 42868 75572
rect 42812 75518 42814 75570
rect 42814 75518 42866 75570
rect 42866 75518 42868 75570
rect 42812 75516 42868 75518
rect 42924 75068 42980 75124
rect 43260 76076 43316 76132
rect 43372 76300 43428 76356
rect 43260 75404 43316 75460
rect 42924 74172 42980 74228
rect 43036 74114 43092 74116
rect 43036 74062 43038 74114
rect 43038 74062 43090 74114
rect 43090 74062 43092 74114
rect 43036 74060 43092 74062
rect 42700 73948 42756 74004
rect 42476 72604 42532 72660
rect 42588 72492 42644 72548
rect 43260 73612 43316 73668
rect 43148 73164 43204 73220
rect 42812 73106 42868 73108
rect 42812 73054 42814 73106
rect 42814 73054 42866 73106
rect 42866 73054 42868 73106
rect 42812 73052 42868 73054
rect 43036 72380 43092 72436
rect 42252 71708 42308 71764
rect 42364 71932 42420 71988
rect 42140 71036 42196 71092
rect 42924 71708 42980 71764
rect 43596 75852 43652 75908
rect 43596 75068 43652 75124
rect 43484 73500 43540 73556
rect 44604 76636 44660 76692
rect 45052 76636 45108 76692
rect 44716 76412 44772 76468
rect 44268 76354 44324 76356
rect 44268 76302 44270 76354
rect 44270 76302 44322 76354
rect 44322 76302 44324 76354
rect 44268 76300 44324 76302
rect 44268 75740 44324 75796
rect 44156 75628 44212 75684
rect 44044 75458 44100 75460
rect 44044 75406 44046 75458
rect 44046 75406 44098 75458
rect 44098 75406 44100 75458
rect 44044 75404 44100 75406
rect 43932 74620 43988 74676
rect 44380 75180 44436 75236
rect 44268 75122 44324 75124
rect 44268 75070 44270 75122
rect 44270 75070 44322 75122
rect 44322 75070 44324 75122
rect 44268 75068 44324 75070
rect 44716 75122 44772 75124
rect 44716 75070 44718 75122
rect 44718 75070 44770 75122
rect 44770 75070 44772 75122
rect 44716 75068 44772 75070
rect 44828 76188 44884 76244
rect 44044 74226 44100 74228
rect 44044 74174 44046 74226
rect 44046 74174 44098 74226
rect 44098 74174 44100 74226
rect 44044 74172 44100 74174
rect 43932 74114 43988 74116
rect 43932 74062 43934 74114
rect 43934 74062 43986 74114
rect 43986 74062 43988 74114
rect 43932 74060 43988 74062
rect 44492 74898 44548 74900
rect 44492 74846 44494 74898
rect 44494 74846 44546 74898
rect 44546 74846 44548 74898
rect 44492 74844 44548 74846
rect 44380 74396 44436 74452
rect 44268 74338 44324 74340
rect 44268 74286 44270 74338
rect 44270 74286 44322 74338
rect 44322 74286 44324 74338
rect 44268 74284 44324 74286
rect 44716 74284 44772 74340
rect 44492 74060 44548 74116
rect 44380 73948 44436 74004
rect 43820 73554 43876 73556
rect 43820 73502 43822 73554
rect 43822 73502 43874 73554
rect 43874 73502 43876 73554
rect 43820 73500 43876 73502
rect 43596 73052 43652 73108
rect 43596 71986 43652 71988
rect 43596 71934 43598 71986
rect 43598 71934 43650 71986
rect 43650 71934 43652 71986
rect 43596 71932 43652 71934
rect 44268 73164 44324 73220
rect 44044 72546 44100 72548
rect 44044 72494 44046 72546
rect 44046 72494 44098 72546
rect 44098 72494 44100 72546
rect 44044 72492 44100 72494
rect 43708 72044 43764 72100
rect 43372 70588 43428 70644
rect 43820 71932 43876 71988
rect 44156 72268 44212 72324
rect 43820 71036 43876 71092
rect 44604 73836 44660 73892
rect 44604 72940 44660 72996
rect 44940 74396 44996 74452
rect 44492 72546 44548 72548
rect 44492 72494 44494 72546
rect 44494 72494 44546 72546
rect 44546 72494 44548 72546
rect 44492 72492 44548 72494
rect 44492 71036 44548 71092
rect 44716 71036 44772 71092
rect 44940 72492 44996 72548
rect 44940 71708 44996 71764
rect 45276 76578 45332 76580
rect 45276 76526 45278 76578
rect 45278 76526 45330 76578
rect 45330 76526 45332 76578
rect 45276 76524 45332 76526
rect 45164 75404 45220 75460
rect 47180 77420 47236 77476
rect 46844 76524 46900 76580
rect 45836 76188 45892 76244
rect 45500 75292 45556 75348
rect 45836 75068 45892 75124
rect 45500 75010 45556 75012
rect 45500 74958 45502 75010
rect 45502 74958 45554 75010
rect 45554 74958 45556 75010
rect 45500 74956 45556 74958
rect 45500 74284 45556 74340
rect 45276 73500 45332 73556
rect 45388 73442 45444 73444
rect 45388 73390 45390 73442
rect 45390 73390 45442 73442
rect 45442 73390 45444 73442
rect 45388 73388 45444 73390
rect 45276 73330 45332 73332
rect 45276 73278 45278 73330
rect 45278 73278 45330 73330
rect 45330 73278 45332 73330
rect 45276 73276 45332 73278
rect 45724 74338 45780 74340
rect 45724 74286 45726 74338
rect 45726 74286 45778 74338
rect 45778 74286 45780 74338
rect 45724 74284 45780 74286
rect 45948 73500 46004 73556
rect 45836 73388 45892 73444
rect 45500 72268 45556 72324
rect 45948 73218 46004 73220
rect 45948 73166 45950 73218
rect 45950 73166 46002 73218
rect 46002 73166 46004 73218
rect 45948 73164 46004 73166
rect 46284 76188 46340 76244
rect 46844 76300 46900 76356
rect 46396 74114 46452 74116
rect 46396 74062 46398 74114
rect 46398 74062 46450 74114
rect 46450 74062 46452 74114
rect 46396 74060 46452 74062
rect 46396 73836 46452 73892
rect 47068 76690 47124 76692
rect 47068 76638 47070 76690
rect 47070 76638 47122 76690
rect 47122 76638 47124 76690
rect 47068 76636 47124 76638
rect 47068 75516 47124 75572
rect 46844 75180 46900 75236
rect 46732 75122 46788 75124
rect 46732 75070 46734 75122
rect 46734 75070 46786 75122
rect 46786 75070 46788 75122
rect 46732 75068 46788 75070
rect 47180 75068 47236 75124
rect 46508 73388 46564 73444
rect 46732 73836 46788 73892
rect 46396 73330 46452 73332
rect 46396 73278 46398 73330
rect 46398 73278 46450 73330
rect 46450 73278 46452 73330
rect 46396 73276 46452 73278
rect 45724 72156 45780 72212
rect 45948 72156 46004 72212
rect 45836 72044 45892 72100
rect 44828 70252 44884 70308
rect 45388 71090 45444 71092
rect 45388 71038 45390 71090
rect 45390 71038 45442 71090
rect 45442 71038 45444 71090
rect 45388 71036 45444 71038
rect 46172 72156 46228 72212
rect 45948 71090 46004 71092
rect 45948 71038 45950 71090
rect 45950 71038 46002 71090
rect 46002 71038 46004 71090
rect 45948 71036 46004 71038
rect 47068 73724 47124 73780
rect 47068 73500 47124 73556
rect 46844 72156 46900 72212
rect 47516 75964 47572 76020
rect 47516 74620 47572 74676
rect 47852 76188 47908 76244
rect 47740 74060 47796 74116
rect 47852 74396 47908 74452
rect 47740 73612 47796 73668
rect 45500 70476 45556 70532
rect 46396 70476 46452 70532
rect 47292 72156 47348 72212
rect 47740 72156 47796 72212
rect 47852 70924 47908 70980
rect 47852 70476 47908 70532
rect 46284 70252 46340 70308
rect 45164 69468 45220 69524
rect 46172 70140 46228 70196
rect 48188 75516 48244 75572
rect 49308 76972 49364 77028
rect 50652 77084 50708 77140
rect 48972 76578 49028 76580
rect 48972 76526 48974 76578
rect 48974 76526 49026 76578
rect 49026 76526 49028 76578
rect 48972 76524 49028 76526
rect 49084 76466 49140 76468
rect 49084 76414 49086 76466
rect 49086 76414 49138 76466
rect 49138 76414 49140 76466
rect 49084 76412 49140 76414
rect 48972 76242 49028 76244
rect 48972 76190 48974 76242
rect 48974 76190 49026 76242
rect 49026 76190 49028 76242
rect 48972 76188 49028 76190
rect 48860 75570 48916 75572
rect 48860 75518 48862 75570
rect 48862 75518 48914 75570
rect 48914 75518 48916 75570
rect 48860 75516 48916 75518
rect 49084 75404 49140 75460
rect 48412 75180 48468 75236
rect 48636 75010 48692 75012
rect 48636 74958 48638 75010
rect 48638 74958 48690 75010
rect 48690 74958 48692 75010
rect 48636 74956 48692 74958
rect 48524 74898 48580 74900
rect 48524 74846 48526 74898
rect 48526 74846 48578 74898
rect 48578 74846 48580 74898
rect 48524 74844 48580 74846
rect 48524 74396 48580 74452
rect 49196 74844 49252 74900
rect 48748 73442 48804 73444
rect 48748 73390 48750 73442
rect 48750 73390 48802 73442
rect 48802 73390 48804 73442
rect 48748 73388 48804 73390
rect 48636 73218 48692 73220
rect 48636 73166 48638 73218
rect 48638 73166 48690 73218
rect 48690 73166 48692 73218
rect 48636 73164 48692 73166
rect 48524 72268 48580 72324
rect 48636 72380 48692 72436
rect 49868 76578 49924 76580
rect 49868 76526 49870 76578
rect 49870 76526 49922 76578
rect 49922 76526 49924 76578
rect 49868 76524 49924 76526
rect 49644 76466 49700 76468
rect 49644 76414 49646 76466
rect 49646 76414 49698 76466
rect 49698 76414 49700 76466
rect 49644 76412 49700 76414
rect 49644 75740 49700 75796
rect 49756 76188 49812 76244
rect 49868 75852 49924 75908
rect 49532 74732 49588 74788
rect 50092 75516 50148 75572
rect 50092 74844 50148 74900
rect 50316 75010 50372 75012
rect 50316 74958 50318 75010
rect 50318 74958 50370 75010
rect 50370 74958 50372 75010
rect 50316 74956 50372 74958
rect 50556 76858 50612 76860
rect 50556 76806 50558 76858
rect 50558 76806 50610 76858
rect 50610 76806 50612 76858
rect 50556 76804 50612 76806
rect 50660 76858 50716 76860
rect 50660 76806 50662 76858
rect 50662 76806 50714 76858
rect 50714 76806 50716 76858
rect 50660 76804 50716 76806
rect 50764 76858 50820 76860
rect 50764 76806 50766 76858
rect 50766 76806 50818 76858
rect 50818 76806 50820 76858
rect 50764 76804 50820 76806
rect 50764 76578 50820 76580
rect 50764 76526 50766 76578
rect 50766 76526 50818 76578
rect 50818 76526 50820 76578
rect 50764 76524 50820 76526
rect 50988 76300 51044 76356
rect 50876 75794 50932 75796
rect 50876 75742 50878 75794
rect 50878 75742 50930 75794
rect 50930 75742 50932 75794
rect 50876 75740 50932 75742
rect 50764 75682 50820 75684
rect 50764 75630 50766 75682
rect 50766 75630 50818 75682
rect 50818 75630 50820 75682
rect 50764 75628 50820 75630
rect 50556 75290 50612 75292
rect 50556 75238 50558 75290
rect 50558 75238 50610 75290
rect 50610 75238 50612 75290
rect 50556 75236 50612 75238
rect 50660 75290 50716 75292
rect 50660 75238 50662 75290
rect 50662 75238 50714 75290
rect 50714 75238 50716 75290
rect 50660 75236 50716 75238
rect 50764 75290 50820 75292
rect 50764 75238 50766 75290
rect 50766 75238 50818 75290
rect 50818 75238 50820 75290
rect 50764 75236 50820 75238
rect 49532 74172 49588 74228
rect 49420 73276 49476 73332
rect 49420 72380 49476 72436
rect 50764 74732 50820 74788
rect 50540 74172 50596 74228
rect 50204 74060 50260 74116
rect 49644 73218 49700 73220
rect 49644 73166 49646 73218
rect 49646 73166 49698 73218
rect 49698 73166 49700 73218
rect 49644 73164 49700 73166
rect 49980 73164 50036 73220
rect 49868 72940 49924 72996
rect 50092 73106 50148 73108
rect 50092 73054 50094 73106
rect 50094 73054 50146 73106
rect 50146 73054 50148 73106
rect 50092 73052 50148 73054
rect 50316 74002 50372 74004
rect 50316 73950 50318 74002
rect 50318 73950 50370 74002
rect 50370 73950 50372 74002
rect 50316 73948 50372 73950
rect 50764 73836 50820 73892
rect 50556 73722 50612 73724
rect 50556 73670 50558 73722
rect 50558 73670 50610 73722
rect 50610 73670 50612 73722
rect 50556 73668 50612 73670
rect 50660 73722 50716 73724
rect 50660 73670 50662 73722
rect 50662 73670 50714 73722
rect 50714 73670 50716 73722
rect 50660 73668 50716 73670
rect 50764 73722 50820 73724
rect 50764 73670 50766 73722
rect 50766 73670 50818 73722
rect 50818 73670 50820 73722
rect 50764 73668 50820 73670
rect 50428 73052 50484 73108
rect 51100 74956 51156 75012
rect 50988 74732 51044 74788
rect 51660 76690 51716 76692
rect 51660 76638 51662 76690
rect 51662 76638 51714 76690
rect 51714 76638 51716 76690
rect 51660 76636 51716 76638
rect 51772 76300 51828 76356
rect 51436 75628 51492 75684
rect 51548 75458 51604 75460
rect 51548 75406 51550 75458
rect 51550 75406 51602 75458
rect 51602 75406 51604 75458
rect 51548 75404 51604 75406
rect 51660 75180 51716 75236
rect 51772 75068 51828 75124
rect 51212 74284 51268 74340
rect 51100 74114 51156 74116
rect 51100 74062 51102 74114
rect 51102 74062 51154 74114
rect 51154 74062 51156 74114
rect 51100 74060 51156 74062
rect 50988 73388 51044 73444
rect 51324 74002 51380 74004
rect 51324 73950 51326 74002
rect 51326 73950 51378 74002
rect 51378 73950 51380 74002
rect 51324 73948 51380 73950
rect 50988 73106 51044 73108
rect 50988 73054 50990 73106
rect 50990 73054 51042 73106
rect 51042 73054 51044 73106
rect 50988 73052 51044 73054
rect 50876 72322 50932 72324
rect 50876 72270 50878 72322
rect 50878 72270 50930 72322
rect 50930 72270 50932 72322
rect 50876 72268 50932 72270
rect 50556 72154 50612 72156
rect 50556 72102 50558 72154
rect 50558 72102 50610 72154
rect 50610 72102 50612 72154
rect 50556 72100 50612 72102
rect 50660 72154 50716 72156
rect 50660 72102 50662 72154
rect 50662 72102 50714 72154
rect 50714 72102 50716 72154
rect 50660 72100 50716 72102
rect 50764 72154 50820 72156
rect 50764 72102 50766 72154
rect 50766 72102 50818 72154
rect 50818 72102 50820 72154
rect 50764 72100 50820 72102
rect 50316 71762 50372 71764
rect 50316 71710 50318 71762
rect 50318 71710 50370 71762
rect 50370 71710 50372 71762
rect 50316 71708 50372 71710
rect 49532 71260 49588 71316
rect 49756 71090 49812 71092
rect 49756 71038 49758 71090
rect 49758 71038 49810 71090
rect 49810 71038 49812 71090
rect 49756 71036 49812 71038
rect 48748 70978 48804 70980
rect 48748 70926 48750 70978
rect 48750 70926 48802 70978
rect 48802 70926 48804 70978
rect 48748 70924 48804 70926
rect 50876 71090 50932 71092
rect 50876 71038 50878 71090
rect 50878 71038 50930 71090
rect 50930 71038 50932 71090
rect 50876 71036 50932 71038
rect 50556 70586 50612 70588
rect 50556 70534 50558 70586
rect 50558 70534 50610 70586
rect 50610 70534 50612 70586
rect 50556 70532 50612 70534
rect 50660 70586 50716 70588
rect 50660 70534 50662 70586
rect 50662 70534 50714 70586
rect 50714 70534 50716 70586
rect 50660 70532 50716 70534
rect 50764 70586 50820 70588
rect 50764 70534 50766 70586
rect 50766 70534 50818 70586
rect 50818 70534 50820 70586
rect 50764 70532 50820 70534
rect 47180 70140 47236 70196
rect 46620 69522 46676 69524
rect 46620 69470 46622 69522
rect 46622 69470 46674 69522
rect 46674 69470 46676 69522
rect 46620 69468 46676 69470
rect 51324 72268 51380 72324
rect 52108 76412 52164 76468
rect 51996 76076 52052 76132
rect 52668 76412 52724 76468
rect 52780 77308 52836 77364
rect 52668 76242 52724 76244
rect 52668 76190 52670 76242
rect 52670 76190 52722 76242
rect 52722 76190 52724 76242
rect 52668 76188 52724 76190
rect 52556 76076 52612 76132
rect 51996 75068 52052 75124
rect 51884 74508 51940 74564
rect 51548 73890 51604 73892
rect 51548 73838 51550 73890
rect 51550 73838 51602 73890
rect 51602 73838 51604 73890
rect 51548 73836 51604 73838
rect 51324 70476 51380 70532
rect 51772 74002 51828 74004
rect 51772 73950 51774 74002
rect 51774 73950 51826 74002
rect 51826 73950 51828 74002
rect 51772 73948 51828 73950
rect 51772 73442 51828 73444
rect 51772 73390 51774 73442
rect 51774 73390 51826 73442
rect 51826 73390 51828 73442
rect 51772 73388 51828 73390
rect 52220 74284 52276 74340
rect 52108 72940 52164 72996
rect 52108 72546 52164 72548
rect 52108 72494 52110 72546
rect 52110 72494 52162 72546
rect 52162 72494 52164 72546
rect 52108 72492 52164 72494
rect 51884 72268 51940 72324
rect 52220 70476 52276 70532
rect 51772 70418 51828 70420
rect 51772 70366 51774 70418
rect 51774 70366 51826 70418
rect 51826 70366 51828 70418
rect 51772 70364 51828 70366
rect 50988 69468 51044 69524
rect 52444 75404 52500 75460
rect 53228 75068 53284 75124
rect 53676 75628 53732 75684
rect 54236 77532 54292 77588
rect 54124 75794 54180 75796
rect 54124 75742 54126 75794
rect 54126 75742 54178 75794
rect 54178 75742 54180 75794
rect 54124 75740 54180 75742
rect 54012 75516 54068 75572
rect 53004 74844 53060 74900
rect 53564 74844 53620 74900
rect 52780 74396 52836 74452
rect 52556 74114 52612 74116
rect 52556 74062 52558 74114
rect 52558 74062 52610 74114
rect 52610 74062 52612 74114
rect 52556 74060 52612 74062
rect 52444 73890 52500 73892
rect 52444 73838 52446 73890
rect 52446 73838 52498 73890
rect 52498 73838 52500 73890
rect 52444 73836 52500 73838
rect 52444 73500 52500 73556
rect 52444 73276 52500 73332
rect 52556 72492 52612 72548
rect 53564 74002 53620 74004
rect 53564 73950 53566 74002
rect 53566 73950 53618 74002
rect 53618 73950 53620 74002
rect 53564 73948 53620 73950
rect 53116 73500 53172 73556
rect 52780 72492 52836 72548
rect 52892 71932 52948 71988
rect 52556 71762 52612 71764
rect 52556 71710 52558 71762
rect 52558 71710 52610 71762
rect 52610 71710 52612 71762
rect 52556 71708 52612 71710
rect 52668 70418 52724 70420
rect 52668 70366 52670 70418
rect 52670 70366 52722 70418
rect 52722 70366 52724 70418
rect 52668 70364 52724 70366
rect 53564 73330 53620 73332
rect 53564 73278 53566 73330
rect 53566 73278 53618 73330
rect 53618 73278 53620 73330
rect 53564 73276 53620 73278
rect 53452 72546 53508 72548
rect 53452 72494 53454 72546
rect 53454 72494 53506 72546
rect 53506 72494 53508 72546
rect 53452 72492 53508 72494
rect 53564 70418 53620 70420
rect 53564 70366 53566 70418
rect 53566 70366 53618 70418
rect 53618 70366 53620 70418
rect 53564 70364 53620 70366
rect 53900 75068 53956 75124
rect 54796 77084 54852 77140
rect 55356 76636 55412 76692
rect 55804 76972 55860 77028
rect 56028 76972 56084 77028
rect 57372 76748 57428 76804
rect 57596 77644 57652 77700
rect 56700 76524 56756 76580
rect 56364 75852 56420 75908
rect 55916 75628 55972 75684
rect 54348 75180 54404 75236
rect 54124 75010 54180 75012
rect 54124 74958 54126 75010
rect 54126 74958 54178 75010
rect 54178 74958 54180 75010
rect 54124 74956 54180 74958
rect 54348 74956 54404 75012
rect 54572 74844 54628 74900
rect 54684 74284 54740 74340
rect 53900 73052 53956 73108
rect 54460 73052 54516 73108
rect 54348 72658 54404 72660
rect 54348 72606 54350 72658
rect 54350 72606 54402 72658
rect 54402 72606 54404 72658
rect 54348 72604 54404 72606
rect 53900 71986 53956 71988
rect 53900 71934 53902 71986
rect 53902 71934 53954 71986
rect 53954 71934 53956 71986
rect 53900 71932 53956 71934
rect 54796 73948 54852 74004
rect 54908 73106 54964 73108
rect 54908 73054 54910 73106
rect 54910 73054 54962 73106
rect 54962 73054 54964 73106
rect 54908 73052 54964 73054
rect 55356 75180 55412 75236
rect 55244 75010 55300 75012
rect 55244 74958 55246 75010
rect 55246 74958 55298 75010
rect 55298 74958 55300 75010
rect 55244 74956 55300 74958
rect 55468 74898 55524 74900
rect 55468 74846 55470 74898
rect 55470 74846 55522 74898
rect 55522 74846 55524 74898
rect 55468 74844 55524 74846
rect 56140 75404 56196 75460
rect 56028 74844 56084 74900
rect 55468 74114 55524 74116
rect 55468 74062 55470 74114
rect 55470 74062 55522 74114
rect 55522 74062 55524 74114
rect 55468 74060 55524 74062
rect 55468 73612 55524 73668
rect 55804 73052 55860 73108
rect 55804 72716 55860 72772
rect 55356 72546 55412 72548
rect 55356 72494 55358 72546
rect 55358 72494 55410 72546
rect 55410 72494 55412 72546
rect 55356 72492 55412 72494
rect 55356 72156 55412 72212
rect 54124 70476 54180 70532
rect 56364 75010 56420 75012
rect 56364 74958 56366 75010
rect 56366 74958 56418 75010
rect 56418 74958 56420 75010
rect 56364 74956 56420 74958
rect 56700 75010 56756 75012
rect 56700 74958 56702 75010
rect 56702 74958 56754 75010
rect 56754 74958 56756 75010
rect 56700 74956 56756 74958
rect 56364 74396 56420 74452
rect 56028 73948 56084 74004
rect 56252 73836 56308 73892
rect 56140 73554 56196 73556
rect 56140 73502 56142 73554
rect 56142 73502 56194 73554
rect 56194 73502 56196 73554
rect 56140 73500 56196 73502
rect 56028 72492 56084 72548
rect 55916 72156 55972 72212
rect 56252 71538 56308 71540
rect 56252 71486 56254 71538
rect 56254 71486 56306 71538
rect 56306 71486 56308 71538
rect 56252 71484 56308 71486
rect 55692 71090 55748 71092
rect 55692 71038 55694 71090
rect 55694 71038 55746 71090
rect 55746 71038 55748 71090
rect 55692 71036 55748 71038
rect 55356 70924 55412 70980
rect 53788 70252 53844 70308
rect 57260 75906 57316 75908
rect 57260 75854 57262 75906
rect 57262 75854 57314 75906
rect 57314 75854 57316 75906
rect 57260 75852 57316 75854
rect 56924 75794 56980 75796
rect 56924 75742 56926 75794
rect 56926 75742 56978 75794
rect 56978 75742 56980 75794
rect 56924 75740 56980 75742
rect 57036 75458 57092 75460
rect 57036 75406 57038 75458
rect 57038 75406 57090 75458
rect 57090 75406 57092 75458
rect 57036 75404 57092 75406
rect 57932 76578 57988 76580
rect 57932 76526 57934 76578
rect 57934 76526 57986 76578
rect 57986 76526 57988 76578
rect 57932 76524 57988 76526
rect 57260 74172 57316 74228
rect 57596 73836 57652 73892
rect 57148 73276 57204 73332
rect 56700 72940 56756 72996
rect 57036 72546 57092 72548
rect 57036 72494 57038 72546
rect 57038 72494 57090 72546
rect 57090 72494 57092 72546
rect 57036 72492 57092 72494
rect 56924 71036 56980 71092
rect 58716 76524 58772 76580
rect 58044 75180 58100 75236
rect 58156 75292 58212 75348
rect 57932 74674 57988 74676
rect 57932 74622 57934 74674
rect 57934 74622 57986 74674
rect 57986 74622 57988 74674
rect 57932 74620 57988 74622
rect 57932 74002 57988 74004
rect 57932 73950 57934 74002
rect 57934 73950 57986 74002
rect 57986 73950 57988 74002
rect 57932 73948 57988 73950
rect 58268 74002 58324 74004
rect 58268 73950 58270 74002
rect 58270 73950 58322 74002
rect 58322 73950 58324 74002
rect 58268 73948 58324 73950
rect 58044 73890 58100 73892
rect 58044 73838 58046 73890
rect 58046 73838 58098 73890
rect 58098 73838 58100 73890
rect 58044 73836 58100 73838
rect 57820 73442 57876 73444
rect 57820 73390 57822 73442
rect 57822 73390 57874 73442
rect 57874 73390 57876 73442
rect 57820 73388 57876 73390
rect 58268 73388 58324 73444
rect 58716 75292 58772 75348
rect 58380 73276 58436 73332
rect 58604 72604 58660 72660
rect 59276 76578 59332 76580
rect 59276 76526 59278 76578
rect 59278 76526 59330 76578
rect 59330 76526 59332 76578
rect 59276 76524 59332 76526
rect 59276 75740 59332 75796
rect 58828 72716 58884 72772
rect 58940 75292 58996 75348
rect 59052 74508 59108 74564
rect 59164 74114 59220 74116
rect 59164 74062 59166 74114
rect 59166 74062 59218 74114
rect 59218 74062 59220 74114
rect 59164 74060 59220 74062
rect 59724 76354 59780 76356
rect 59724 76302 59726 76354
rect 59726 76302 59778 76354
rect 59778 76302 59780 76354
rect 59724 76300 59780 76302
rect 59948 75740 60004 75796
rect 59612 75458 59668 75460
rect 59612 75406 59614 75458
rect 59614 75406 59666 75458
rect 59666 75406 59668 75458
rect 59612 75404 59668 75406
rect 59388 74508 59444 74564
rect 59052 72604 59108 72660
rect 59500 73388 59556 73444
rect 59388 72940 59444 72996
rect 59836 74508 59892 74564
rect 59724 73836 59780 73892
rect 59836 74060 59892 74116
rect 60508 75570 60564 75572
rect 60508 75518 60510 75570
rect 60510 75518 60562 75570
rect 60562 75518 60564 75570
rect 60508 75516 60564 75518
rect 60284 74620 60340 74676
rect 60732 75010 60788 75012
rect 60732 74958 60734 75010
rect 60734 74958 60786 75010
rect 60786 74958 60788 75010
rect 60732 74956 60788 74958
rect 60060 73724 60116 73780
rect 60284 73442 60340 73444
rect 60284 73390 60286 73442
rect 60286 73390 60338 73442
rect 60338 73390 60340 73442
rect 60284 73388 60340 73390
rect 60620 74002 60676 74004
rect 60620 73950 60622 74002
rect 60622 73950 60674 74002
rect 60674 73950 60676 74002
rect 60620 73948 60676 73950
rect 60732 73612 60788 73668
rect 60844 73724 60900 73780
rect 60508 73500 60564 73556
rect 60956 73500 61012 73556
rect 61068 74508 61124 74564
rect 59276 72546 59332 72548
rect 59276 72494 59278 72546
rect 59278 72494 59330 72546
rect 59330 72494 59332 72546
rect 59276 72492 59332 72494
rect 58268 71484 58324 71540
rect 58940 71090 58996 71092
rect 58940 71038 58942 71090
rect 58942 71038 58994 71090
rect 58994 71038 58996 71090
rect 58940 71036 58996 71038
rect 60284 72658 60340 72660
rect 60284 72606 60286 72658
rect 60286 72606 60338 72658
rect 60338 72606 60340 72658
rect 60284 72604 60340 72606
rect 59836 71036 59892 71092
rect 61292 75682 61348 75684
rect 61292 75630 61294 75682
rect 61294 75630 61346 75682
rect 61346 75630 61348 75682
rect 61292 75628 61348 75630
rect 61852 76690 61908 76692
rect 61852 76638 61854 76690
rect 61854 76638 61906 76690
rect 61906 76638 61908 76690
rect 61852 76636 61908 76638
rect 61852 76188 61908 76244
rect 61628 75852 61684 75908
rect 61404 75068 61460 75124
rect 61516 75458 61572 75460
rect 61516 75406 61518 75458
rect 61518 75406 61570 75458
rect 61570 75406 61572 75458
rect 61516 75404 61572 75406
rect 61180 74284 61236 74340
rect 61292 74172 61348 74228
rect 62524 76972 62580 77028
rect 62076 75516 62132 75572
rect 61964 75180 62020 75236
rect 62412 75628 62468 75684
rect 62188 74956 62244 75012
rect 62300 74620 62356 74676
rect 61852 74396 61908 74452
rect 61852 73948 61908 74004
rect 61404 73890 61460 73892
rect 61404 73838 61406 73890
rect 61406 73838 61458 73890
rect 61458 73838 61460 73890
rect 61404 73836 61460 73838
rect 61404 73554 61460 73556
rect 61404 73502 61406 73554
rect 61406 73502 61458 73554
rect 61458 73502 61460 73554
rect 61404 73500 61460 73502
rect 63196 76748 63252 76804
rect 62860 75794 62916 75796
rect 62860 75742 62862 75794
rect 62862 75742 62914 75794
rect 62914 75742 62916 75794
rect 62860 75740 62916 75742
rect 62748 75292 62804 75348
rect 62636 75122 62692 75124
rect 62636 75070 62638 75122
rect 62638 75070 62690 75122
rect 62690 75070 62692 75122
rect 62636 75068 62692 75070
rect 62300 73554 62356 73556
rect 62300 73502 62302 73554
rect 62302 73502 62354 73554
rect 62354 73502 62356 73554
rect 62300 73500 62356 73502
rect 63308 75516 63364 75572
rect 63756 76466 63812 76468
rect 63756 76414 63758 76466
rect 63758 76414 63810 76466
rect 63810 76414 63812 76466
rect 63756 76412 63812 76414
rect 64428 76578 64484 76580
rect 64428 76526 64430 76578
rect 64430 76526 64482 76578
rect 64482 76526 64484 76578
rect 64428 76524 64484 76526
rect 64764 76524 64820 76580
rect 64764 75740 64820 75796
rect 64092 75404 64148 75460
rect 63420 75068 63476 75124
rect 63980 75122 64036 75124
rect 63980 75070 63982 75122
rect 63982 75070 64034 75122
rect 64034 75070 64036 75122
rect 63980 75068 64036 75070
rect 62860 74620 62916 74676
rect 64540 74620 64596 74676
rect 63308 74284 63364 74340
rect 65324 75740 65380 75796
rect 64988 75292 65044 75348
rect 65916 76074 65972 76076
rect 65916 76022 65918 76074
rect 65918 76022 65970 76074
rect 65970 76022 65972 76074
rect 65916 76020 65972 76022
rect 66020 76074 66076 76076
rect 66020 76022 66022 76074
rect 66022 76022 66074 76074
rect 66074 76022 66076 76074
rect 66020 76020 66076 76022
rect 66124 76074 66180 76076
rect 66124 76022 66126 76074
rect 66126 76022 66178 76074
rect 66178 76022 66180 76074
rect 66124 76020 66180 76022
rect 65436 75516 65492 75572
rect 65996 75458 66052 75460
rect 65996 75406 65998 75458
rect 65998 75406 66050 75458
rect 66050 75406 66052 75458
rect 65996 75404 66052 75406
rect 67228 76578 67284 76580
rect 67228 76526 67230 76578
rect 67230 76526 67282 76578
rect 67282 76526 67284 76578
rect 67228 76524 67284 76526
rect 66780 75740 66836 75796
rect 66668 75570 66724 75572
rect 66668 75518 66670 75570
rect 66670 75518 66722 75570
rect 66722 75518 66724 75570
rect 66668 75516 66724 75518
rect 67452 75516 67508 75572
rect 68012 75570 68068 75572
rect 68012 75518 68014 75570
rect 68014 75518 68066 75570
rect 68066 75518 68068 75570
rect 68012 75516 68068 75518
rect 66332 75404 66388 75460
rect 67340 75458 67396 75460
rect 67340 75406 67342 75458
rect 67342 75406 67394 75458
rect 67394 75406 67396 75458
rect 67340 75404 67396 75406
rect 68348 76242 68404 76244
rect 68348 76190 68350 76242
rect 68350 76190 68402 76242
rect 68402 76190 68404 76242
rect 68348 76188 68404 76190
rect 68684 75794 68740 75796
rect 68684 75742 68686 75794
rect 68686 75742 68738 75794
rect 68738 75742 68740 75794
rect 68684 75740 68740 75742
rect 69356 76300 69412 76356
rect 70140 76524 70196 76580
rect 70588 75740 70644 75796
rect 69468 75516 69524 75572
rect 70252 75570 70308 75572
rect 70252 75518 70254 75570
rect 70254 75518 70306 75570
rect 70306 75518 70308 75570
rect 70252 75516 70308 75518
rect 70924 77420 70980 77476
rect 72156 76860 72212 76916
rect 71484 76748 71540 76804
rect 72380 76748 72436 76804
rect 71484 76578 71540 76580
rect 71484 76526 71486 76578
rect 71486 76526 71538 76578
rect 71538 76526 71540 76578
rect 71484 76524 71540 76526
rect 73052 77308 73108 77364
rect 73500 76636 73556 76692
rect 73948 76860 74004 76916
rect 74620 76690 74676 76692
rect 74620 76638 74622 76690
rect 74622 76638 74674 76690
rect 74674 76638 74676 76690
rect 74620 76636 74676 76638
rect 70812 75516 70868 75572
rect 68796 75404 68852 75460
rect 69132 75404 69188 75460
rect 69692 75458 69748 75460
rect 69692 75406 69694 75458
rect 69694 75406 69746 75458
rect 69746 75406 69748 75458
rect 69692 75404 69748 75406
rect 73052 75570 73108 75572
rect 73052 75518 73054 75570
rect 73054 75518 73106 75570
rect 73106 75518 73108 75570
rect 73052 75516 73108 75518
rect 73948 75682 74004 75684
rect 73948 75630 73950 75682
rect 73950 75630 74002 75682
rect 74002 75630 74004 75682
rect 73948 75628 74004 75630
rect 75516 76636 75572 76692
rect 76300 76690 76356 76692
rect 76300 76638 76302 76690
rect 76302 76638 76354 76690
rect 76354 76638 76356 76690
rect 76300 76636 76356 76638
rect 74844 75516 74900 75572
rect 76076 75570 76132 75572
rect 76076 75518 76078 75570
rect 76078 75518 76130 75570
rect 76130 75518 76132 75570
rect 76076 75516 76132 75518
rect 77196 75570 77252 75572
rect 77196 75518 77198 75570
rect 77198 75518 77250 75570
rect 77250 75518 77252 75570
rect 77196 75516 77252 75518
rect 76860 74956 76916 75012
rect 77644 75010 77700 75012
rect 77644 74958 77646 75010
rect 77646 74958 77698 75010
rect 77698 74958 77700 75010
rect 77644 74956 77700 74958
rect 78092 74956 78148 75012
rect 74508 74674 74564 74676
rect 74508 74622 74510 74674
rect 74510 74622 74562 74674
rect 74562 74622 74564 74674
rect 74508 74620 74564 74622
rect 65916 74506 65972 74508
rect 65916 74454 65918 74506
rect 65918 74454 65970 74506
rect 65970 74454 65972 74506
rect 65916 74452 65972 74454
rect 66020 74506 66076 74508
rect 66020 74454 66022 74506
rect 66022 74454 66074 74506
rect 66074 74454 66076 74506
rect 66020 74452 66076 74454
rect 66124 74506 66180 74508
rect 66124 74454 66126 74506
rect 66126 74454 66178 74506
rect 66178 74454 66180 74506
rect 66124 74452 66180 74454
rect 64876 73948 64932 74004
rect 65916 72938 65972 72940
rect 65916 72886 65918 72938
rect 65918 72886 65970 72938
rect 65970 72886 65972 72938
rect 65916 72884 65972 72886
rect 66020 72938 66076 72940
rect 66020 72886 66022 72938
rect 66022 72886 66074 72938
rect 66074 72886 66076 72938
rect 66020 72884 66076 72886
rect 66124 72938 66180 72940
rect 66124 72886 66126 72938
rect 66126 72886 66178 72938
rect 66178 72886 66180 72938
rect 66124 72884 66180 72886
rect 61964 72604 62020 72660
rect 65916 71370 65972 71372
rect 65916 71318 65918 71370
rect 65918 71318 65970 71370
rect 65970 71318 65972 71370
rect 65916 71316 65972 71318
rect 66020 71370 66076 71372
rect 66020 71318 66022 71370
rect 66022 71318 66074 71370
rect 66074 71318 66076 71370
rect 66020 71316 66076 71318
rect 66124 71370 66180 71372
rect 66124 71318 66126 71370
rect 66126 71318 66178 71370
rect 66178 71318 66180 71370
rect 66124 71316 66180 71318
rect 60508 70476 60564 70532
rect 65916 69802 65972 69804
rect 65916 69750 65918 69802
rect 65918 69750 65970 69802
rect 65970 69750 65972 69802
rect 65916 69748 65972 69750
rect 66020 69802 66076 69804
rect 66020 69750 66022 69802
rect 66022 69750 66074 69802
rect 66074 69750 66076 69802
rect 66020 69748 66076 69750
rect 66124 69802 66180 69804
rect 66124 69750 66126 69802
rect 66126 69750 66178 69802
rect 66178 69750 66180 69802
rect 66124 69748 66180 69750
rect 52780 69522 52836 69524
rect 52780 69470 52782 69522
rect 52782 69470 52834 69522
rect 52834 69470 52836 69522
rect 52780 69468 52836 69470
rect 19836 69018 19892 69020
rect 19836 68966 19838 69018
rect 19838 68966 19890 69018
rect 19890 68966 19892 69018
rect 19836 68964 19892 68966
rect 19940 69018 19996 69020
rect 19940 68966 19942 69018
rect 19942 68966 19994 69018
rect 19994 68966 19996 69018
rect 19940 68964 19996 68966
rect 20044 69018 20100 69020
rect 20044 68966 20046 69018
rect 20046 68966 20098 69018
rect 20098 68966 20100 69018
rect 20044 68964 20100 68966
rect 50556 69018 50612 69020
rect 50556 68966 50558 69018
rect 50558 68966 50610 69018
rect 50610 68966 50612 69018
rect 50556 68964 50612 68966
rect 50660 69018 50716 69020
rect 50660 68966 50662 69018
rect 50662 68966 50714 69018
rect 50714 68966 50716 69018
rect 50660 68964 50716 68966
rect 50764 69018 50820 69020
rect 50764 68966 50766 69018
rect 50766 68966 50818 69018
rect 50818 68966 50820 69018
rect 50764 68964 50820 68966
rect 4476 68234 4532 68236
rect 4476 68182 4478 68234
rect 4478 68182 4530 68234
rect 4530 68182 4532 68234
rect 4476 68180 4532 68182
rect 4580 68234 4636 68236
rect 4580 68182 4582 68234
rect 4582 68182 4634 68234
rect 4634 68182 4636 68234
rect 4580 68180 4636 68182
rect 4684 68234 4740 68236
rect 4684 68182 4686 68234
rect 4686 68182 4738 68234
rect 4738 68182 4740 68234
rect 4684 68180 4740 68182
rect 35196 68234 35252 68236
rect 35196 68182 35198 68234
rect 35198 68182 35250 68234
rect 35250 68182 35252 68234
rect 35196 68180 35252 68182
rect 35300 68234 35356 68236
rect 35300 68182 35302 68234
rect 35302 68182 35354 68234
rect 35354 68182 35356 68234
rect 35300 68180 35356 68182
rect 35404 68234 35460 68236
rect 35404 68182 35406 68234
rect 35406 68182 35458 68234
rect 35458 68182 35460 68234
rect 35404 68180 35460 68182
rect 65916 68234 65972 68236
rect 65916 68182 65918 68234
rect 65918 68182 65970 68234
rect 65970 68182 65972 68234
rect 65916 68180 65972 68182
rect 66020 68234 66076 68236
rect 66020 68182 66022 68234
rect 66022 68182 66074 68234
rect 66074 68182 66076 68234
rect 66020 68180 66076 68182
rect 66124 68234 66180 68236
rect 66124 68182 66126 68234
rect 66126 68182 66178 68234
rect 66178 68182 66180 68234
rect 66124 68180 66180 68182
rect 19836 67450 19892 67452
rect 19836 67398 19838 67450
rect 19838 67398 19890 67450
rect 19890 67398 19892 67450
rect 19836 67396 19892 67398
rect 19940 67450 19996 67452
rect 19940 67398 19942 67450
rect 19942 67398 19994 67450
rect 19994 67398 19996 67450
rect 19940 67396 19996 67398
rect 20044 67450 20100 67452
rect 20044 67398 20046 67450
rect 20046 67398 20098 67450
rect 20098 67398 20100 67450
rect 20044 67396 20100 67398
rect 50556 67450 50612 67452
rect 50556 67398 50558 67450
rect 50558 67398 50610 67450
rect 50610 67398 50612 67450
rect 50556 67396 50612 67398
rect 50660 67450 50716 67452
rect 50660 67398 50662 67450
rect 50662 67398 50714 67450
rect 50714 67398 50716 67450
rect 50660 67396 50716 67398
rect 50764 67450 50820 67452
rect 50764 67398 50766 67450
rect 50766 67398 50818 67450
rect 50818 67398 50820 67450
rect 50764 67396 50820 67398
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 35196 66666 35252 66668
rect 35196 66614 35198 66666
rect 35198 66614 35250 66666
rect 35250 66614 35252 66666
rect 35196 66612 35252 66614
rect 35300 66666 35356 66668
rect 35300 66614 35302 66666
rect 35302 66614 35354 66666
rect 35354 66614 35356 66666
rect 35300 66612 35356 66614
rect 35404 66666 35460 66668
rect 35404 66614 35406 66666
rect 35406 66614 35458 66666
rect 35458 66614 35460 66666
rect 35404 66612 35460 66614
rect 65916 66666 65972 66668
rect 65916 66614 65918 66666
rect 65918 66614 65970 66666
rect 65970 66614 65972 66666
rect 65916 66612 65972 66614
rect 66020 66666 66076 66668
rect 66020 66614 66022 66666
rect 66022 66614 66074 66666
rect 66074 66614 66076 66666
rect 66020 66612 66076 66614
rect 66124 66666 66180 66668
rect 66124 66614 66126 66666
rect 66126 66614 66178 66666
rect 66178 66614 66180 66666
rect 66124 66612 66180 66614
rect 19836 65882 19892 65884
rect 19836 65830 19838 65882
rect 19838 65830 19890 65882
rect 19890 65830 19892 65882
rect 19836 65828 19892 65830
rect 19940 65882 19996 65884
rect 19940 65830 19942 65882
rect 19942 65830 19994 65882
rect 19994 65830 19996 65882
rect 19940 65828 19996 65830
rect 20044 65882 20100 65884
rect 20044 65830 20046 65882
rect 20046 65830 20098 65882
rect 20098 65830 20100 65882
rect 20044 65828 20100 65830
rect 50556 65882 50612 65884
rect 50556 65830 50558 65882
rect 50558 65830 50610 65882
rect 50610 65830 50612 65882
rect 50556 65828 50612 65830
rect 50660 65882 50716 65884
rect 50660 65830 50662 65882
rect 50662 65830 50714 65882
rect 50714 65830 50716 65882
rect 50660 65828 50716 65830
rect 50764 65882 50820 65884
rect 50764 65830 50766 65882
rect 50766 65830 50818 65882
rect 50818 65830 50820 65882
rect 50764 65828 50820 65830
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 35196 65098 35252 65100
rect 35196 65046 35198 65098
rect 35198 65046 35250 65098
rect 35250 65046 35252 65098
rect 35196 65044 35252 65046
rect 35300 65098 35356 65100
rect 35300 65046 35302 65098
rect 35302 65046 35354 65098
rect 35354 65046 35356 65098
rect 35300 65044 35356 65046
rect 35404 65098 35460 65100
rect 35404 65046 35406 65098
rect 35406 65046 35458 65098
rect 35458 65046 35460 65098
rect 35404 65044 35460 65046
rect 65916 65098 65972 65100
rect 65916 65046 65918 65098
rect 65918 65046 65970 65098
rect 65970 65046 65972 65098
rect 65916 65044 65972 65046
rect 66020 65098 66076 65100
rect 66020 65046 66022 65098
rect 66022 65046 66074 65098
rect 66074 65046 66076 65098
rect 66020 65044 66076 65046
rect 66124 65098 66180 65100
rect 66124 65046 66126 65098
rect 66126 65046 66178 65098
rect 66178 65046 66180 65098
rect 66124 65044 66180 65046
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 50556 64314 50612 64316
rect 50556 64262 50558 64314
rect 50558 64262 50610 64314
rect 50610 64262 50612 64314
rect 50556 64260 50612 64262
rect 50660 64314 50716 64316
rect 50660 64262 50662 64314
rect 50662 64262 50714 64314
rect 50714 64262 50716 64314
rect 50660 64260 50716 64262
rect 50764 64314 50820 64316
rect 50764 64262 50766 64314
rect 50766 64262 50818 64314
rect 50818 64262 50820 64314
rect 50764 64260 50820 64262
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 35404 63476 35460 63478
rect 65916 63530 65972 63532
rect 65916 63478 65918 63530
rect 65918 63478 65970 63530
rect 65970 63478 65972 63530
rect 65916 63476 65972 63478
rect 66020 63530 66076 63532
rect 66020 63478 66022 63530
rect 66022 63478 66074 63530
rect 66074 63478 66076 63530
rect 66020 63476 66076 63478
rect 66124 63530 66180 63532
rect 66124 63478 66126 63530
rect 66126 63478 66178 63530
rect 66178 63478 66180 63530
rect 66124 63476 66180 63478
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 50556 62746 50612 62748
rect 50556 62694 50558 62746
rect 50558 62694 50610 62746
rect 50610 62694 50612 62746
rect 50556 62692 50612 62694
rect 50660 62746 50716 62748
rect 50660 62694 50662 62746
rect 50662 62694 50714 62746
rect 50714 62694 50716 62746
rect 50660 62692 50716 62694
rect 50764 62746 50820 62748
rect 50764 62694 50766 62746
rect 50766 62694 50818 62746
rect 50818 62694 50820 62746
rect 50764 62692 50820 62694
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 65916 61962 65972 61964
rect 65916 61910 65918 61962
rect 65918 61910 65970 61962
rect 65970 61910 65972 61962
rect 65916 61908 65972 61910
rect 66020 61962 66076 61964
rect 66020 61910 66022 61962
rect 66022 61910 66074 61962
rect 66074 61910 66076 61962
rect 66020 61908 66076 61910
rect 66124 61962 66180 61964
rect 66124 61910 66126 61962
rect 66126 61910 66178 61962
rect 66178 61910 66180 61962
rect 66124 61908 66180 61910
rect 19836 61178 19892 61180
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 50556 61178 50612 61180
rect 50556 61126 50558 61178
rect 50558 61126 50610 61178
rect 50610 61126 50612 61178
rect 50556 61124 50612 61126
rect 50660 61178 50716 61180
rect 50660 61126 50662 61178
rect 50662 61126 50714 61178
rect 50714 61126 50716 61178
rect 50660 61124 50716 61126
rect 50764 61178 50820 61180
rect 50764 61126 50766 61178
rect 50766 61126 50818 61178
rect 50818 61126 50820 61178
rect 50764 61124 50820 61126
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 65916 60394 65972 60396
rect 65916 60342 65918 60394
rect 65918 60342 65970 60394
rect 65970 60342 65972 60394
rect 65916 60340 65972 60342
rect 66020 60394 66076 60396
rect 66020 60342 66022 60394
rect 66022 60342 66074 60394
rect 66074 60342 66076 60394
rect 66020 60340 66076 60342
rect 66124 60394 66180 60396
rect 66124 60342 66126 60394
rect 66126 60342 66178 60394
rect 66178 60342 66180 60394
rect 66124 60340 66180 60342
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 50556 59610 50612 59612
rect 50556 59558 50558 59610
rect 50558 59558 50610 59610
rect 50610 59558 50612 59610
rect 50556 59556 50612 59558
rect 50660 59610 50716 59612
rect 50660 59558 50662 59610
rect 50662 59558 50714 59610
rect 50714 59558 50716 59610
rect 50660 59556 50716 59558
rect 50764 59610 50820 59612
rect 50764 59558 50766 59610
rect 50766 59558 50818 59610
rect 50818 59558 50820 59610
rect 50764 59556 50820 59558
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 65916 58826 65972 58828
rect 65916 58774 65918 58826
rect 65918 58774 65970 58826
rect 65970 58774 65972 58826
rect 65916 58772 65972 58774
rect 66020 58826 66076 58828
rect 66020 58774 66022 58826
rect 66022 58774 66074 58826
rect 66074 58774 66076 58826
rect 66020 58772 66076 58774
rect 66124 58826 66180 58828
rect 66124 58774 66126 58826
rect 66126 58774 66178 58826
rect 66178 58774 66180 58826
rect 66124 58772 66180 58774
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 50556 58042 50612 58044
rect 50556 57990 50558 58042
rect 50558 57990 50610 58042
rect 50610 57990 50612 58042
rect 50556 57988 50612 57990
rect 50660 58042 50716 58044
rect 50660 57990 50662 58042
rect 50662 57990 50714 58042
rect 50714 57990 50716 58042
rect 50660 57988 50716 57990
rect 50764 58042 50820 58044
rect 50764 57990 50766 58042
rect 50766 57990 50818 58042
rect 50818 57990 50820 58042
rect 50764 57988 50820 57990
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 65916 57258 65972 57260
rect 65916 57206 65918 57258
rect 65918 57206 65970 57258
rect 65970 57206 65972 57258
rect 65916 57204 65972 57206
rect 66020 57258 66076 57260
rect 66020 57206 66022 57258
rect 66022 57206 66074 57258
rect 66074 57206 66076 57258
rect 66020 57204 66076 57206
rect 66124 57258 66180 57260
rect 66124 57206 66126 57258
rect 66126 57206 66178 57258
rect 66178 57206 66180 57258
rect 66124 57204 66180 57206
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 65916 55690 65972 55692
rect 65916 55638 65918 55690
rect 65918 55638 65970 55690
rect 65970 55638 65972 55690
rect 65916 55636 65972 55638
rect 66020 55690 66076 55692
rect 66020 55638 66022 55690
rect 66022 55638 66074 55690
rect 66074 55638 66076 55690
rect 66020 55636 66076 55638
rect 66124 55690 66180 55692
rect 66124 55638 66126 55690
rect 66126 55638 66178 55690
rect 66178 55638 66180 55690
rect 66124 55636 66180 55638
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 65916 54122 65972 54124
rect 65916 54070 65918 54122
rect 65918 54070 65970 54122
rect 65970 54070 65972 54122
rect 65916 54068 65972 54070
rect 66020 54122 66076 54124
rect 66020 54070 66022 54122
rect 66022 54070 66074 54122
rect 66074 54070 66076 54122
rect 66020 54068 66076 54070
rect 66124 54122 66180 54124
rect 66124 54070 66126 54122
rect 66126 54070 66178 54122
rect 66178 54070 66180 54122
rect 66124 54068 66180 54070
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 65916 52554 65972 52556
rect 65916 52502 65918 52554
rect 65918 52502 65970 52554
rect 65970 52502 65972 52554
rect 65916 52500 65972 52502
rect 66020 52554 66076 52556
rect 66020 52502 66022 52554
rect 66022 52502 66074 52554
rect 66074 52502 66076 52554
rect 66020 52500 66076 52502
rect 66124 52554 66180 52556
rect 66124 52502 66126 52554
rect 66126 52502 66178 52554
rect 66178 52502 66180 52554
rect 66124 52500 66180 52502
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 65916 50986 65972 50988
rect 65916 50934 65918 50986
rect 65918 50934 65970 50986
rect 65970 50934 65972 50986
rect 65916 50932 65972 50934
rect 66020 50986 66076 50988
rect 66020 50934 66022 50986
rect 66022 50934 66074 50986
rect 66074 50934 66076 50986
rect 66020 50932 66076 50934
rect 66124 50986 66180 50988
rect 66124 50934 66126 50986
rect 66126 50934 66178 50986
rect 66178 50934 66180 50986
rect 66124 50932 66180 50934
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 65916 49418 65972 49420
rect 65916 49366 65918 49418
rect 65918 49366 65970 49418
rect 65970 49366 65972 49418
rect 65916 49364 65972 49366
rect 66020 49418 66076 49420
rect 66020 49366 66022 49418
rect 66022 49366 66074 49418
rect 66074 49366 66076 49418
rect 66020 49364 66076 49366
rect 66124 49418 66180 49420
rect 66124 49366 66126 49418
rect 66126 49366 66178 49418
rect 66178 49366 66180 49418
rect 66124 49364 66180 49366
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 65916 47850 65972 47852
rect 65916 47798 65918 47850
rect 65918 47798 65970 47850
rect 65970 47798 65972 47850
rect 65916 47796 65972 47798
rect 66020 47850 66076 47852
rect 66020 47798 66022 47850
rect 66022 47798 66074 47850
rect 66074 47798 66076 47850
rect 66020 47796 66076 47798
rect 66124 47850 66180 47852
rect 66124 47798 66126 47850
rect 66126 47798 66178 47850
rect 66178 47798 66180 47850
rect 66124 47796 66180 47798
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 65916 46282 65972 46284
rect 65916 46230 65918 46282
rect 65918 46230 65970 46282
rect 65970 46230 65972 46282
rect 65916 46228 65972 46230
rect 66020 46282 66076 46284
rect 66020 46230 66022 46282
rect 66022 46230 66074 46282
rect 66074 46230 66076 46282
rect 66020 46228 66076 46230
rect 66124 46282 66180 46284
rect 66124 46230 66126 46282
rect 66126 46230 66178 46282
rect 66178 46230 66180 46282
rect 66124 46228 66180 46230
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 65916 44714 65972 44716
rect 65916 44662 65918 44714
rect 65918 44662 65970 44714
rect 65970 44662 65972 44714
rect 65916 44660 65972 44662
rect 66020 44714 66076 44716
rect 66020 44662 66022 44714
rect 66022 44662 66074 44714
rect 66074 44662 66076 44714
rect 66020 44660 66076 44662
rect 66124 44714 66180 44716
rect 66124 44662 66126 44714
rect 66126 44662 66178 44714
rect 66178 44662 66180 44714
rect 66124 44660 66180 44662
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 65916 43146 65972 43148
rect 65916 43094 65918 43146
rect 65918 43094 65970 43146
rect 65970 43094 65972 43146
rect 65916 43092 65972 43094
rect 66020 43146 66076 43148
rect 66020 43094 66022 43146
rect 66022 43094 66074 43146
rect 66074 43094 66076 43146
rect 66020 43092 66076 43094
rect 66124 43146 66180 43148
rect 66124 43094 66126 43146
rect 66126 43094 66178 43146
rect 66178 43094 66180 43146
rect 66124 43092 66180 43094
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 65916 41578 65972 41580
rect 65916 41526 65918 41578
rect 65918 41526 65970 41578
rect 65970 41526 65972 41578
rect 65916 41524 65972 41526
rect 66020 41578 66076 41580
rect 66020 41526 66022 41578
rect 66022 41526 66074 41578
rect 66074 41526 66076 41578
rect 66020 41524 66076 41526
rect 66124 41578 66180 41580
rect 66124 41526 66126 41578
rect 66126 41526 66178 41578
rect 66178 41526 66180 41578
rect 66124 41524 66180 41526
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 65916 40010 65972 40012
rect 65916 39958 65918 40010
rect 65918 39958 65970 40010
rect 65970 39958 65972 40010
rect 65916 39956 65972 39958
rect 66020 40010 66076 40012
rect 66020 39958 66022 40010
rect 66022 39958 66074 40010
rect 66074 39958 66076 40010
rect 66020 39956 66076 39958
rect 66124 40010 66180 40012
rect 66124 39958 66126 40010
rect 66126 39958 66178 40010
rect 66178 39958 66180 40010
rect 66124 39956 66180 39958
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 65916 38442 65972 38444
rect 65916 38390 65918 38442
rect 65918 38390 65970 38442
rect 65970 38390 65972 38442
rect 65916 38388 65972 38390
rect 66020 38442 66076 38444
rect 66020 38390 66022 38442
rect 66022 38390 66074 38442
rect 66074 38390 66076 38442
rect 66020 38388 66076 38390
rect 66124 38442 66180 38444
rect 66124 38390 66126 38442
rect 66126 38390 66178 38442
rect 66178 38390 66180 38442
rect 66124 38388 66180 38390
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 65916 36874 65972 36876
rect 65916 36822 65918 36874
rect 65918 36822 65970 36874
rect 65970 36822 65972 36874
rect 65916 36820 65972 36822
rect 66020 36874 66076 36876
rect 66020 36822 66022 36874
rect 66022 36822 66074 36874
rect 66074 36822 66076 36874
rect 66020 36820 66076 36822
rect 66124 36874 66180 36876
rect 66124 36822 66126 36874
rect 66126 36822 66178 36874
rect 66178 36822 66180 36874
rect 66124 36820 66180 36822
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 65916 35306 65972 35308
rect 65916 35254 65918 35306
rect 65918 35254 65970 35306
rect 65970 35254 65972 35306
rect 65916 35252 65972 35254
rect 66020 35306 66076 35308
rect 66020 35254 66022 35306
rect 66022 35254 66074 35306
rect 66074 35254 66076 35306
rect 66020 35252 66076 35254
rect 66124 35306 66180 35308
rect 66124 35254 66126 35306
rect 66126 35254 66178 35306
rect 66178 35254 66180 35306
rect 66124 35252 66180 35254
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 65916 33738 65972 33740
rect 65916 33686 65918 33738
rect 65918 33686 65970 33738
rect 65970 33686 65972 33738
rect 65916 33684 65972 33686
rect 66020 33738 66076 33740
rect 66020 33686 66022 33738
rect 66022 33686 66074 33738
rect 66074 33686 66076 33738
rect 66020 33684 66076 33686
rect 66124 33738 66180 33740
rect 66124 33686 66126 33738
rect 66126 33686 66178 33738
rect 66178 33686 66180 33738
rect 66124 33684 66180 33686
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 65916 32170 65972 32172
rect 65916 32118 65918 32170
rect 65918 32118 65970 32170
rect 65970 32118 65972 32170
rect 65916 32116 65972 32118
rect 66020 32170 66076 32172
rect 66020 32118 66022 32170
rect 66022 32118 66074 32170
rect 66074 32118 66076 32170
rect 66020 32116 66076 32118
rect 66124 32170 66180 32172
rect 66124 32118 66126 32170
rect 66126 32118 66178 32170
rect 66178 32118 66180 32170
rect 66124 32116 66180 32118
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 65916 30602 65972 30604
rect 65916 30550 65918 30602
rect 65918 30550 65970 30602
rect 65970 30550 65972 30602
rect 65916 30548 65972 30550
rect 66020 30602 66076 30604
rect 66020 30550 66022 30602
rect 66022 30550 66074 30602
rect 66074 30550 66076 30602
rect 66020 30548 66076 30550
rect 66124 30602 66180 30604
rect 66124 30550 66126 30602
rect 66126 30550 66178 30602
rect 66178 30550 66180 30602
rect 66124 30548 66180 30550
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 65916 29034 65972 29036
rect 65916 28982 65918 29034
rect 65918 28982 65970 29034
rect 65970 28982 65972 29034
rect 65916 28980 65972 28982
rect 66020 29034 66076 29036
rect 66020 28982 66022 29034
rect 66022 28982 66074 29034
rect 66074 28982 66076 29034
rect 66020 28980 66076 28982
rect 66124 29034 66180 29036
rect 66124 28982 66126 29034
rect 66126 28982 66178 29034
rect 66178 28982 66180 29034
rect 66124 28980 66180 28982
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 65916 27466 65972 27468
rect 65916 27414 65918 27466
rect 65918 27414 65970 27466
rect 65970 27414 65972 27466
rect 65916 27412 65972 27414
rect 66020 27466 66076 27468
rect 66020 27414 66022 27466
rect 66022 27414 66074 27466
rect 66074 27414 66076 27466
rect 66020 27412 66076 27414
rect 66124 27466 66180 27468
rect 66124 27414 66126 27466
rect 66126 27414 66178 27466
rect 66178 27414 66180 27466
rect 66124 27412 66180 27414
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 65916 25898 65972 25900
rect 65916 25846 65918 25898
rect 65918 25846 65970 25898
rect 65970 25846 65972 25898
rect 65916 25844 65972 25846
rect 66020 25898 66076 25900
rect 66020 25846 66022 25898
rect 66022 25846 66074 25898
rect 66074 25846 66076 25898
rect 66020 25844 66076 25846
rect 66124 25898 66180 25900
rect 66124 25846 66126 25898
rect 66126 25846 66178 25898
rect 66178 25846 66180 25898
rect 66124 25844 66180 25846
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 65916 24330 65972 24332
rect 65916 24278 65918 24330
rect 65918 24278 65970 24330
rect 65970 24278 65972 24330
rect 65916 24276 65972 24278
rect 66020 24330 66076 24332
rect 66020 24278 66022 24330
rect 66022 24278 66074 24330
rect 66074 24278 66076 24330
rect 66020 24276 66076 24278
rect 66124 24330 66180 24332
rect 66124 24278 66126 24330
rect 66126 24278 66178 24330
rect 66178 24278 66180 24330
rect 66124 24276 66180 24278
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 65916 22762 65972 22764
rect 65916 22710 65918 22762
rect 65918 22710 65970 22762
rect 65970 22710 65972 22762
rect 65916 22708 65972 22710
rect 66020 22762 66076 22764
rect 66020 22710 66022 22762
rect 66022 22710 66074 22762
rect 66074 22710 66076 22762
rect 66020 22708 66076 22710
rect 66124 22762 66180 22764
rect 66124 22710 66126 22762
rect 66126 22710 66178 22762
rect 66178 22710 66180 22762
rect 66124 22708 66180 22710
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 65916 21194 65972 21196
rect 65916 21142 65918 21194
rect 65918 21142 65970 21194
rect 65970 21142 65972 21194
rect 65916 21140 65972 21142
rect 66020 21194 66076 21196
rect 66020 21142 66022 21194
rect 66022 21142 66074 21194
rect 66074 21142 66076 21194
rect 66020 21140 66076 21142
rect 66124 21194 66180 21196
rect 66124 21142 66126 21194
rect 66126 21142 66178 21194
rect 66178 21142 66180 21194
rect 66124 21140 66180 21142
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 65916 19626 65972 19628
rect 65916 19574 65918 19626
rect 65918 19574 65970 19626
rect 65970 19574 65972 19626
rect 65916 19572 65972 19574
rect 66020 19626 66076 19628
rect 66020 19574 66022 19626
rect 66022 19574 66074 19626
rect 66074 19574 66076 19626
rect 66020 19572 66076 19574
rect 66124 19626 66180 19628
rect 66124 19574 66126 19626
rect 66126 19574 66178 19626
rect 66178 19574 66180 19626
rect 66124 19572 66180 19574
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 65916 18058 65972 18060
rect 65916 18006 65918 18058
rect 65918 18006 65970 18058
rect 65970 18006 65972 18058
rect 65916 18004 65972 18006
rect 66020 18058 66076 18060
rect 66020 18006 66022 18058
rect 66022 18006 66074 18058
rect 66074 18006 66076 18058
rect 66020 18004 66076 18006
rect 66124 18058 66180 18060
rect 66124 18006 66126 18058
rect 66126 18006 66178 18058
rect 66178 18006 66180 18058
rect 66124 18004 66180 18006
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 65916 16490 65972 16492
rect 65916 16438 65918 16490
rect 65918 16438 65970 16490
rect 65970 16438 65972 16490
rect 65916 16436 65972 16438
rect 66020 16490 66076 16492
rect 66020 16438 66022 16490
rect 66022 16438 66074 16490
rect 66074 16438 66076 16490
rect 66020 16436 66076 16438
rect 66124 16490 66180 16492
rect 66124 16438 66126 16490
rect 66126 16438 66178 16490
rect 66178 16438 66180 16490
rect 66124 16436 66180 16438
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 65916 14922 65972 14924
rect 65916 14870 65918 14922
rect 65918 14870 65970 14922
rect 65970 14870 65972 14922
rect 65916 14868 65972 14870
rect 66020 14922 66076 14924
rect 66020 14870 66022 14922
rect 66022 14870 66074 14922
rect 66074 14870 66076 14922
rect 66020 14868 66076 14870
rect 66124 14922 66180 14924
rect 66124 14870 66126 14922
rect 66126 14870 66178 14922
rect 66178 14870 66180 14922
rect 66124 14868 66180 14870
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 65916 13354 65972 13356
rect 65916 13302 65918 13354
rect 65918 13302 65970 13354
rect 65970 13302 65972 13354
rect 65916 13300 65972 13302
rect 66020 13354 66076 13356
rect 66020 13302 66022 13354
rect 66022 13302 66074 13354
rect 66074 13302 66076 13354
rect 66020 13300 66076 13302
rect 66124 13354 66180 13356
rect 66124 13302 66126 13354
rect 66126 13302 66178 13354
rect 66178 13302 66180 13354
rect 66124 13300 66180 13302
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 65916 11786 65972 11788
rect 65916 11734 65918 11786
rect 65918 11734 65970 11786
rect 65970 11734 65972 11786
rect 65916 11732 65972 11734
rect 66020 11786 66076 11788
rect 66020 11734 66022 11786
rect 66022 11734 66074 11786
rect 66074 11734 66076 11786
rect 66020 11732 66076 11734
rect 66124 11786 66180 11788
rect 66124 11734 66126 11786
rect 66126 11734 66178 11786
rect 66178 11734 66180 11786
rect 66124 11732 66180 11734
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 65916 10218 65972 10220
rect 65916 10166 65918 10218
rect 65918 10166 65970 10218
rect 65970 10166 65972 10218
rect 65916 10164 65972 10166
rect 66020 10218 66076 10220
rect 66020 10166 66022 10218
rect 66022 10166 66074 10218
rect 66074 10166 66076 10218
rect 66020 10164 66076 10166
rect 66124 10218 66180 10220
rect 66124 10166 66126 10218
rect 66126 10166 66178 10218
rect 66178 10166 66180 10218
rect 66124 10164 66180 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 65916 8650 65972 8652
rect 65916 8598 65918 8650
rect 65918 8598 65970 8650
rect 65970 8598 65972 8650
rect 65916 8596 65972 8598
rect 66020 8650 66076 8652
rect 66020 8598 66022 8650
rect 66022 8598 66074 8650
rect 66074 8598 66076 8650
rect 66020 8596 66076 8598
rect 66124 8650 66180 8652
rect 66124 8598 66126 8650
rect 66126 8598 66178 8650
rect 66178 8598 66180 8650
rect 66124 8596 66180 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 65916 7082 65972 7084
rect 65916 7030 65918 7082
rect 65918 7030 65970 7082
rect 65970 7030 65972 7082
rect 65916 7028 65972 7030
rect 66020 7082 66076 7084
rect 66020 7030 66022 7082
rect 66022 7030 66074 7082
rect 66074 7030 66076 7082
rect 66020 7028 66076 7030
rect 66124 7082 66180 7084
rect 66124 7030 66126 7082
rect 66126 7030 66178 7082
rect 66178 7030 66180 7082
rect 66124 7028 66180 7030
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 65916 5514 65972 5516
rect 65916 5462 65918 5514
rect 65918 5462 65970 5514
rect 65970 5462 65972 5514
rect 65916 5460 65972 5462
rect 66020 5514 66076 5516
rect 66020 5462 66022 5514
rect 66022 5462 66074 5514
rect 66074 5462 66076 5514
rect 66020 5460 66076 5462
rect 66124 5514 66180 5516
rect 66124 5462 66126 5514
rect 66126 5462 66178 5514
rect 66178 5462 66180 5514
rect 66124 5460 66180 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 45052 3276 45108 3332
rect 45612 3330 45668 3332
rect 45612 3278 45614 3330
rect 45614 3278 45666 3330
rect 45666 3278 45668 3330
rect 45612 3276 45668 3278
rect 47740 3276 47796 3332
rect 48860 3330 48916 3332
rect 48860 3278 48862 3330
rect 48862 3278 48914 3330
rect 48914 3278 48916 3330
rect 48860 3276 48916 3278
rect 48412 1708 48468 1764
rect 49532 1708 49588 1764
rect 49756 3276 49812 3332
rect 50876 3330 50932 3332
rect 50876 3278 50878 3330
rect 50878 3278 50930 3330
rect 50930 3278 50932 3330
rect 50876 3276 50932 3278
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 51772 3276 51828 3332
rect 52780 3330 52836 3332
rect 52780 3278 52782 3330
rect 52782 3278 52834 3330
rect 52834 3278 52836 3330
rect 52780 3276 52836 3278
rect 53116 3276 53172 3332
rect 54124 3330 54180 3332
rect 54124 3278 54126 3330
rect 54126 3278 54178 3330
rect 54178 3278 54180 3330
rect 54124 3276 54180 3278
rect 54460 3276 54516 3332
rect 55468 3330 55524 3332
rect 55468 3278 55470 3330
rect 55470 3278 55522 3330
rect 55522 3278 55524 3330
rect 55468 3276 55524 3278
rect 56476 3276 56532 3332
rect 57372 3330 57428 3332
rect 57372 3278 57374 3330
rect 57374 3278 57426 3330
rect 57426 3278 57428 3330
rect 57372 3276 57428 3278
rect 58492 3276 58548 3332
rect 59388 3330 59444 3332
rect 59388 3278 59390 3330
rect 59390 3278 59442 3330
rect 59442 3278 59444 3330
rect 59388 3276 59444 3278
rect 59836 3276 59892 3332
rect 60620 3330 60676 3332
rect 60620 3278 60622 3330
rect 60622 3278 60674 3330
rect 60674 3278 60676 3330
rect 60620 3276 60676 3278
rect 61852 3276 61908 3332
rect 62636 3330 62692 3332
rect 62636 3278 62638 3330
rect 62638 3278 62690 3330
rect 62690 3278 62692 3330
rect 62636 3276 62692 3278
rect 65916 3946 65972 3948
rect 65916 3894 65918 3946
rect 65918 3894 65970 3946
rect 65970 3894 65972 3946
rect 65916 3892 65972 3894
rect 66020 3946 66076 3948
rect 66020 3894 66022 3946
rect 66022 3894 66074 3946
rect 66074 3894 66076 3946
rect 66020 3892 66076 3894
rect 66124 3946 66180 3948
rect 66124 3894 66126 3946
rect 66126 3894 66178 3946
rect 66178 3894 66180 3946
rect 66124 3892 66180 3894
rect 65324 3276 65380 3332
rect 65884 3330 65940 3332
rect 65884 3278 65886 3330
rect 65886 3278 65938 3330
rect 65938 3278 65940 3330
rect 65884 3276 65940 3278
rect 66668 3276 66724 3332
rect 67228 3330 67284 3332
rect 67228 3278 67230 3330
rect 67230 3278 67282 3330
rect 67282 3278 67284 3330
rect 67228 3276 67284 3278
rect 67900 3276 67956 3332
rect 69132 3330 69188 3332
rect 69132 3278 69134 3330
rect 69134 3278 69186 3330
rect 69186 3278 69188 3330
rect 69132 3276 69188 3278
rect 68572 1708 68628 1764
rect 69804 1708 69860 1764
rect 69916 1820 69972 1876
rect 71148 1820 71204 1876
rect 71260 3276 71316 3332
rect 72380 3330 72436 3332
rect 72380 3278 72382 3330
rect 72382 3278 72434 3330
rect 72434 3278 72436 3330
rect 72380 3276 72436 3278
rect 71932 1708 71988 1764
rect 73052 1708 73108 1764
rect 73500 4396 73556 4452
rect 73276 3276 73332 3332
rect 74060 4450 74116 4452
rect 74060 4398 74062 4450
rect 74062 4398 74114 4450
rect 74114 4398 74116 4450
rect 74060 4396 74116 4398
rect 74396 3330 74452 3332
rect 74396 3278 74398 3330
rect 74398 3278 74450 3330
rect 74450 3278 74452 3330
rect 74396 3276 74452 3278
<< metal3 >>
rect 34402 77644 34412 77700
rect 34468 77644 57596 77700
rect 57652 77644 57662 77700
rect 35634 77532 35644 77588
rect 35700 77532 54236 77588
rect 54292 77532 54302 77588
rect 47170 77420 47180 77476
rect 47236 77420 70924 77476
rect 70980 77420 70990 77476
rect 52770 77308 52780 77364
rect 52836 77308 73052 77364
rect 73108 77308 73118 77364
rect 50642 77084 50652 77140
rect 50708 77084 54796 77140
rect 54852 77084 54862 77140
rect 49298 76972 49308 77028
rect 49364 76972 55804 77028
rect 55860 76972 55870 77028
rect 56018 76972 56028 77028
rect 56084 76972 62524 77028
rect 62580 76972 62590 77028
rect 72146 76860 72156 76916
rect 72212 76860 73948 76916
rect 74004 76860 74014 76916
rect 19826 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20110 76860
rect 50546 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50830 76860
rect 57362 76748 57372 76804
rect 57428 76748 63196 76804
rect 63252 76748 63262 76804
rect 71474 76748 71484 76804
rect 71540 76748 72380 76804
rect 72436 76748 72446 76804
rect 2930 76636 2940 76692
rect 2996 76636 3836 76692
rect 3892 76636 3902 76692
rect 6850 76636 6860 76692
rect 6916 76636 7980 76692
rect 8036 76636 43372 76692
rect 43428 76636 43438 76692
rect 44594 76636 44604 76692
rect 44660 76636 45052 76692
rect 45108 76636 47068 76692
rect 47124 76636 47134 76692
rect 47292 76636 51660 76692
rect 51716 76636 51726 76692
rect 55346 76636 55356 76692
rect 55412 76636 61852 76692
rect 61908 76636 61918 76692
rect 73490 76636 73500 76692
rect 73556 76636 74620 76692
rect 74676 76636 74686 76692
rect 75506 76636 75516 76692
rect 75572 76636 76300 76692
rect 76356 76636 76366 76692
rect 47292 76580 47348 76636
rect 3602 76524 3612 76580
rect 3668 76524 5852 76580
rect 5908 76524 5918 76580
rect 38546 76524 38556 76580
rect 38612 76524 38892 76580
rect 38948 76524 38958 76580
rect 39228 76524 40404 76580
rect 40562 76524 40572 76580
rect 40628 76524 41132 76580
rect 41188 76524 42028 76580
rect 42084 76524 42094 76580
rect 42578 76524 42588 76580
rect 42644 76524 45276 76580
rect 45332 76524 45342 76580
rect 46834 76524 46844 76580
rect 46900 76524 47348 76580
rect 48962 76524 48972 76580
rect 49028 76524 49868 76580
rect 49924 76524 50764 76580
rect 50820 76524 50830 76580
rect 56690 76524 56700 76580
rect 56756 76524 57932 76580
rect 57988 76524 57998 76580
rect 58706 76524 58716 76580
rect 58772 76524 59276 76580
rect 59332 76524 64428 76580
rect 64484 76524 64494 76580
rect 64754 76524 64764 76580
rect 64820 76524 67228 76580
rect 67284 76524 67294 76580
rect 70130 76524 70140 76580
rect 70196 76524 71484 76580
rect 71540 76524 71550 76580
rect 39228 76468 39284 76524
rect 40348 76468 40404 76524
rect 14914 76412 14924 76468
rect 14980 76412 15820 76468
rect 15876 76412 15886 76468
rect 18834 76412 18844 76468
rect 18900 76412 19852 76468
rect 19908 76412 19918 76468
rect 37202 76412 37212 76468
rect 37268 76412 39284 76468
rect 39340 76412 40124 76468
rect 40180 76412 40190 76468
rect 40348 76412 41692 76468
rect 41748 76412 41758 76468
rect 39340 76356 39396 76412
rect 42812 76356 42868 76524
rect 57932 76468 57988 76524
rect 43026 76412 43036 76468
rect 43092 76412 44716 76468
rect 44772 76412 44782 76468
rect 49074 76412 49084 76468
rect 49140 76412 49644 76468
rect 49700 76412 49710 76468
rect 52098 76412 52108 76468
rect 52164 76412 52668 76468
rect 52724 76412 52734 76468
rect 57932 76412 63756 76468
rect 63812 76412 63822 76468
rect 37090 76300 37100 76356
rect 37156 76300 37884 76356
rect 37940 76300 39396 76356
rect 39554 76300 39564 76356
rect 39620 76300 41020 76356
rect 41076 76300 41086 76356
rect 42812 76300 43372 76356
rect 43428 76300 43438 76356
rect 44258 76300 44268 76356
rect 44324 76300 46844 76356
rect 46900 76300 46910 76356
rect 50978 76300 50988 76356
rect 51044 76300 51772 76356
rect 51828 76300 59724 76356
rect 59780 76300 69356 76356
rect 69412 76300 69422 76356
rect 19842 76188 19852 76244
rect 19908 76188 34300 76244
rect 34356 76188 34366 76244
rect 37202 76188 37212 76244
rect 37268 76188 39452 76244
rect 39508 76188 39518 76244
rect 40338 76188 40348 76244
rect 40404 76188 41468 76244
rect 41524 76188 41534 76244
rect 41682 76188 41692 76244
rect 41748 76188 44828 76244
rect 44884 76188 45836 76244
rect 45892 76188 46284 76244
rect 46340 76188 46350 76244
rect 47842 76188 47852 76244
rect 47908 76188 48972 76244
rect 49028 76188 49038 76244
rect 49746 76188 49756 76244
rect 49812 76188 52668 76244
rect 52724 76188 52734 76244
rect 61842 76188 61852 76244
rect 61908 76188 68348 76244
rect 68404 76188 68414 76244
rect 42466 76076 42476 76132
rect 42532 76076 43260 76132
rect 43316 76076 51996 76132
rect 52052 76076 52556 76132
rect 52612 76076 52622 76132
rect 4466 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4750 76076
rect 35186 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35470 76076
rect 65906 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66190 76076
rect 20850 75964 20860 76020
rect 20916 75964 34188 76020
rect 34244 75964 34254 76020
rect 36082 75964 36092 76020
rect 36148 75964 47516 76020
rect 47572 75964 47582 76020
rect 3378 75852 3388 75908
rect 3444 75852 21756 75908
rect 21812 75852 21822 75908
rect 22754 75852 22764 75908
rect 22820 75852 23996 75908
rect 24052 75852 36204 75908
rect 36260 75852 36270 75908
rect 43586 75852 43596 75908
rect 43652 75852 49868 75908
rect 49924 75852 49934 75908
rect 56354 75852 56364 75908
rect 56420 75852 57260 75908
rect 57316 75852 61628 75908
rect 61684 75852 61694 75908
rect 24770 75740 24780 75796
rect 24836 75740 28476 75796
rect 28532 75740 28542 75796
rect 29138 75740 29148 75796
rect 29204 75740 29214 75796
rect 31826 75740 31836 75796
rect 31892 75740 32732 75796
rect 32788 75740 32798 75796
rect 39442 75740 39452 75796
rect 39508 75740 40012 75796
rect 40068 75740 40078 75796
rect 41682 75740 41692 75796
rect 41748 75740 44268 75796
rect 44324 75740 44334 75796
rect 49634 75740 49644 75796
rect 49700 75740 50876 75796
rect 50932 75740 50942 75796
rect 54114 75740 54124 75796
rect 54180 75740 56924 75796
rect 56980 75740 56990 75796
rect 59266 75740 59276 75796
rect 59332 75740 59948 75796
rect 60004 75740 62860 75796
rect 62916 75740 62926 75796
rect 64754 75740 64764 75796
rect 64820 75740 65324 75796
rect 65380 75740 65390 75796
rect 66770 75740 66780 75796
rect 66836 75740 68684 75796
rect 68740 75740 70588 75796
rect 70644 75740 70654 75796
rect 16706 75628 16716 75684
rect 16772 75628 17836 75684
rect 17892 75628 23492 75684
rect 13010 75516 13020 75572
rect 13076 75516 13692 75572
rect 13748 75516 13758 75572
rect 21074 75516 21084 75572
rect 21140 75516 21644 75572
rect 21700 75516 21710 75572
rect 15810 75404 15820 75460
rect 15876 75404 21420 75460
rect 21476 75404 21486 75460
rect 19826 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20110 75292
rect 23436 75236 23492 75628
rect 29148 75572 29204 75740
rect 30034 75628 30044 75684
rect 30100 75628 30940 75684
rect 30996 75628 31006 75684
rect 37660 75628 39620 75684
rect 39778 75628 39788 75684
rect 39844 75628 40684 75684
rect 40740 75628 40750 75684
rect 43026 75628 43036 75684
rect 43092 75628 44156 75684
rect 44212 75628 44222 75684
rect 50754 75628 50764 75684
rect 50820 75628 51436 75684
rect 51492 75628 51502 75684
rect 53666 75628 53676 75684
rect 53732 75628 55916 75684
rect 55972 75628 61292 75684
rect 61348 75628 61358 75684
rect 62402 75628 62412 75684
rect 62468 75628 73948 75684
rect 74004 75628 74014 75684
rect 27906 75516 27916 75572
rect 27972 75516 29204 75572
rect 29922 75516 29932 75572
rect 29988 75516 33180 75572
rect 33236 75516 33246 75572
rect 37660 75460 37716 75628
rect 39564 75572 39620 75628
rect 39564 75516 40796 75572
rect 40852 75516 40862 75572
rect 41794 75516 41804 75572
rect 41860 75516 41870 75572
rect 42242 75516 42252 75572
rect 42308 75516 42812 75572
rect 42868 75516 42878 75572
rect 47058 75516 47068 75572
rect 47124 75516 48188 75572
rect 48244 75516 48860 75572
rect 48916 75516 48926 75572
rect 50082 75516 50092 75572
rect 50148 75516 52724 75572
rect 54002 75516 54012 75572
rect 54068 75516 60508 75572
rect 60564 75516 60574 75572
rect 62066 75516 62076 75572
rect 62132 75516 63308 75572
rect 63364 75516 63374 75572
rect 65426 75516 65436 75572
rect 65492 75516 66668 75572
rect 66724 75516 66734 75572
rect 67442 75516 67452 75572
rect 67508 75516 68012 75572
rect 68068 75516 68078 75572
rect 69458 75516 69468 75572
rect 69524 75516 70252 75572
rect 70308 75516 70318 75572
rect 70802 75516 70812 75572
rect 70868 75516 73052 75572
rect 73108 75516 73118 75572
rect 74834 75516 74844 75572
rect 74900 75516 76076 75572
rect 76132 75516 77196 75572
rect 77252 75516 77262 75572
rect 41804 75460 41860 75516
rect 52668 75460 52724 75516
rect 28130 75404 28140 75460
rect 28196 75404 30156 75460
rect 30212 75404 30222 75460
rect 30482 75404 30492 75460
rect 30548 75404 31500 75460
rect 31556 75404 32844 75460
rect 32900 75404 32910 75460
rect 37650 75404 37660 75460
rect 37716 75404 37726 75460
rect 40226 75404 40236 75460
rect 40292 75404 43260 75460
rect 43316 75404 44044 75460
rect 44100 75404 44110 75460
rect 45154 75404 45164 75460
rect 45220 75404 49084 75460
rect 49140 75404 49150 75460
rect 51538 75404 51548 75460
rect 51604 75404 52444 75460
rect 52500 75404 52510 75460
rect 52668 75404 55468 75460
rect 56130 75404 56140 75460
rect 56196 75404 57036 75460
rect 57092 75404 59612 75460
rect 59668 75404 61516 75460
rect 61572 75404 61582 75460
rect 64082 75404 64092 75460
rect 64148 75404 65996 75460
rect 66052 75404 66062 75460
rect 66322 75404 66332 75460
rect 66388 75404 67340 75460
rect 67396 75404 67406 75460
rect 68786 75404 68796 75460
rect 68852 75404 69132 75460
rect 69188 75404 69692 75460
rect 69748 75404 69758 75460
rect 30156 75348 30212 75404
rect 55412 75348 55468 75404
rect 30156 75292 30716 75348
rect 30772 75292 30782 75348
rect 39666 75292 39676 75348
rect 39732 75292 45500 75348
rect 45556 75292 45566 75348
rect 55412 75292 58156 75348
rect 58212 75292 58716 75348
rect 58772 75292 58940 75348
rect 58996 75292 59006 75348
rect 62738 75292 62748 75348
rect 62804 75292 64988 75348
rect 65044 75292 65054 75348
rect 50546 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50830 75292
rect 23436 75180 30940 75236
rect 30996 75180 31006 75236
rect 31154 75180 31164 75236
rect 31220 75180 40124 75236
rect 40180 75180 40190 75236
rect 44370 75180 44380 75236
rect 44436 75180 46844 75236
rect 46900 75180 48412 75236
rect 48468 75180 48478 75236
rect 51622 75180 51660 75236
rect 51716 75180 51726 75236
rect 54338 75180 54348 75236
rect 54404 75180 55356 75236
rect 55412 75180 55422 75236
rect 58034 75180 58044 75236
rect 58100 75180 61964 75236
rect 62020 75180 62030 75236
rect 30258 75068 30268 75124
rect 30324 75068 31500 75124
rect 31556 75068 32060 75124
rect 32116 75068 32126 75124
rect 33058 75068 33068 75124
rect 33124 75068 34412 75124
rect 34468 75068 34478 75124
rect 35746 75068 35756 75124
rect 35812 75068 39900 75124
rect 39956 75068 39966 75124
rect 42914 75068 42924 75124
rect 42980 75068 43596 75124
rect 43652 75068 44268 75124
rect 44324 75068 44334 75124
rect 44594 75068 44604 75124
rect 44660 75068 44716 75124
rect 44772 75068 44782 75124
rect 45826 75068 45836 75124
rect 45892 75068 46732 75124
rect 46788 75068 47180 75124
rect 47236 75068 47246 75124
rect 51762 75068 51772 75124
rect 51828 75068 51996 75124
rect 52052 75068 52062 75124
rect 53218 75068 53228 75124
rect 53284 75068 53900 75124
rect 53956 75068 54404 75124
rect 61394 75068 61404 75124
rect 61460 75068 62636 75124
rect 62692 75068 62702 75124
rect 63410 75068 63420 75124
rect 63476 75068 63980 75124
rect 64036 75068 64046 75124
rect 54348 75012 54404 75068
rect 33730 74956 33740 75012
rect 33796 74956 37940 75012
rect 38770 74956 38780 75012
rect 38836 74956 40572 75012
rect 40628 74956 40638 75012
rect 40786 74956 40796 75012
rect 40852 74956 45500 75012
rect 45556 74956 45566 75012
rect 48626 74956 48636 75012
rect 48692 74956 50316 75012
rect 50372 74956 50382 75012
rect 51090 74956 51100 75012
rect 51156 74956 54124 75012
rect 54180 74956 54190 75012
rect 54338 74956 54348 75012
rect 54404 74956 55244 75012
rect 55300 74956 56364 75012
rect 56420 74956 56430 75012
rect 56690 74956 56700 75012
rect 56756 74956 60732 75012
rect 60788 74956 62188 75012
rect 62244 74956 62254 75012
rect 76850 74956 76860 75012
rect 76916 74956 77644 75012
rect 77700 74956 78092 75012
rect 78148 74956 78158 75012
rect 37884 74900 37940 74956
rect 54124 74900 54180 74956
rect 30706 74844 30716 74900
rect 30772 74844 32060 74900
rect 32116 74844 32126 74900
rect 34514 74844 34524 74900
rect 34580 74844 35644 74900
rect 35700 74844 35710 74900
rect 36082 74844 36092 74900
rect 36148 74844 36988 74900
rect 37044 74844 37054 74900
rect 37874 74844 37884 74900
rect 37940 74844 38444 74900
rect 38500 74844 38892 74900
rect 38948 74844 39676 74900
rect 39732 74844 39742 74900
rect 41654 74844 41692 74900
rect 41748 74844 41758 74900
rect 42354 74844 42364 74900
rect 42420 74844 44492 74900
rect 44548 74844 44558 74900
rect 48514 74844 48524 74900
rect 48580 74844 49196 74900
rect 49252 74844 50092 74900
rect 50148 74844 50158 74900
rect 52994 74844 53004 74900
rect 53060 74844 53564 74900
rect 53620 74844 53630 74900
rect 54124 74844 54572 74900
rect 54628 74844 54638 74900
rect 55458 74844 55468 74900
rect 55524 74844 56028 74900
rect 56084 74844 56094 74900
rect 32610 74732 32620 74788
rect 32676 74732 34076 74788
rect 34132 74732 36428 74788
rect 36484 74732 36494 74788
rect 49522 74732 49532 74788
rect 49588 74732 50764 74788
rect 50820 74732 50830 74788
rect 50978 74732 50988 74788
rect 51044 74732 51940 74788
rect 43922 74620 43932 74676
rect 43988 74620 47516 74676
rect 47572 74620 47582 74676
rect 51884 74564 51940 74732
rect 57922 74620 57932 74676
rect 57988 74620 60284 74676
rect 60340 74620 60350 74676
rect 62290 74620 62300 74676
rect 62356 74620 62860 74676
rect 62916 74620 64540 74676
rect 64596 74620 74508 74676
rect 74564 74620 74574 74676
rect 62300 74564 62356 74620
rect 36754 74508 36764 74564
rect 36820 74508 36988 74564
rect 37044 74508 37996 74564
rect 38052 74508 38062 74564
rect 51874 74508 51884 74564
rect 51940 74508 51950 74564
rect 59042 74508 59052 74564
rect 59108 74508 59388 74564
rect 59444 74508 59836 74564
rect 59892 74508 61068 74564
rect 61124 74508 62356 74564
rect 4466 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4750 74508
rect 35186 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35470 74508
rect 65906 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66190 74508
rect 26562 74396 26572 74452
rect 26628 74396 31948 74452
rect 32004 74396 32620 74452
rect 32676 74396 32686 74452
rect 35634 74396 35644 74452
rect 35700 74396 42140 74452
rect 42196 74396 42206 74452
rect 44370 74396 44380 74452
rect 44436 74396 44940 74452
rect 44996 74396 45006 74452
rect 45724 74396 47852 74452
rect 47908 74396 48524 74452
rect 48580 74396 52780 74452
rect 52836 74396 52846 74452
rect 56354 74396 56364 74452
rect 56420 74396 61852 74452
rect 61908 74396 61918 74452
rect 45724 74340 45780 74396
rect 56364 74340 56420 74396
rect 21746 74284 21756 74340
rect 21812 74284 28812 74340
rect 28868 74284 28878 74340
rect 29362 74284 29372 74340
rect 29428 74284 34188 74340
rect 34244 74284 34254 74340
rect 36530 74284 36540 74340
rect 36596 74284 40684 74340
rect 40740 74284 40750 74340
rect 42242 74284 42252 74340
rect 42308 74284 44268 74340
rect 44324 74284 44716 74340
rect 44772 74284 44782 74340
rect 45490 74284 45500 74340
rect 45556 74284 45724 74340
rect 45780 74284 45790 74340
rect 51202 74284 51212 74340
rect 51268 74284 51660 74340
rect 51716 74284 51726 74340
rect 52182 74284 52220 74340
rect 52276 74284 52286 74340
rect 54674 74284 54684 74340
rect 54740 74284 56420 74340
rect 61170 74284 61180 74340
rect 61236 74284 63308 74340
rect 63364 74284 63374 74340
rect 28578 74172 28588 74228
rect 28644 74172 29708 74228
rect 29764 74172 31164 74228
rect 31220 74172 31230 74228
rect 32162 74172 32172 74228
rect 32228 74172 33852 74228
rect 33908 74172 33918 74228
rect 34290 74172 34300 74228
rect 34356 74172 34524 74228
rect 34580 74172 35308 74228
rect 35364 74172 35374 74228
rect 40114 74172 40124 74228
rect 40180 74172 40852 74228
rect 40796 74116 40852 74172
rect 41804 74172 42924 74228
rect 42980 74172 44044 74228
rect 44100 74172 44110 74228
rect 45836 74172 49532 74228
rect 49588 74172 49598 74228
rect 50530 74172 50540 74228
rect 50596 74172 51828 74228
rect 57250 74172 57260 74228
rect 57316 74172 61292 74228
rect 61348 74172 61358 74228
rect 34738 74060 34748 74116
rect 34804 74060 35980 74116
rect 36036 74060 37548 74116
rect 37604 74060 37614 74116
rect 37762 74060 37772 74116
rect 37828 74060 38108 74116
rect 38164 74060 40460 74116
rect 40516 74060 40526 74116
rect 40786 74060 40796 74116
rect 40852 74060 41580 74116
rect 41636 74060 41646 74116
rect 41804 74004 41860 74172
rect 45836 74116 45892 74172
rect 43026 74060 43036 74116
rect 43092 74060 43932 74116
rect 43988 74060 43998 74116
rect 44482 74060 44492 74116
rect 44548 74060 45836 74116
rect 45892 74060 45902 74116
rect 46386 74060 46396 74116
rect 46452 74060 47740 74116
rect 47796 74060 47806 74116
rect 50194 74060 50204 74116
rect 50260 74060 51100 74116
rect 51156 74060 51166 74116
rect 51772 74004 51828 74172
rect 52546 74060 52556 74116
rect 52612 74060 55468 74116
rect 55524 74060 55534 74116
rect 59154 74060 59164 74116
rect 59220 74060 59836 74116
rect 59892 74060 61908 74116
rect 61852 74004 61908 74060
rect 28802 73948 28812 74004
rect 28868 73948 29484 74004
rect 29540 73948 30156 74004
rect 30212 73948 31052 74004
rect 31108 73948 31118 74004
rect 34626 73948 34636 74004
rect 34692 73948 35420 74004
rect 35476 73948 35486 74004
rect 36876 73948 39004 74004
rect 39060 73948 39070 74004
rect 40562 73948 40572 74004
rect 40628 73948 41804 74004
rect 41860 73948 41870 74004
rect 42690 73948 42700 74004
rect 42756 73948 44380 74004
rect 44436 73948 44446 74004
rect 50306 73948 50316 74004
rect 50372 73948 51324 74004
rect 51380 73948 51390 74004
rect 51762 73948 51772 74004
rect 51828 73948 53564 74004
rect 53620 73948 54796 74004
rect 54852 73948 54862 74004
rect 56018 73948 56028 74004
rect 56084 73948 57932 74004
rect 57988 73948 57998 74004
rect 58258 73948 58268 74004
rect 58324 73948 60620 74004
rect 60676 73948 60686 74004
rect 61842 73948 61852 74004
rect 61908 73948 64876 74004
rect 64932 73948 64942 74004
rect 36876 73892 36932 73948
rect 31378 73836 31388 73892
rect 31444 73836 33292 73892
rect 33348 73836 33358 73892
rect 36866 73836 36876 73892
rect 36932 73836 36942 73892
rect 44594 73836 44604 73892
rect 44660 73836 46396 73892
rect 46452 73836 46732 73892
rect 46788 73836 46798 73892
rect 50754 73836 50764 73892
rect 50820 73836 51548 73892
rect 51604 73836 51614 73892
rect 52210 73836 52220 73892
rect 52276 73836 52444 73892
rect 52500 73836 52510 73892
rect 56242 73836 56252 73892
rect 56308 73836 57596 73892
rect 57652 73836 58044 73892
rect 58100 73836 58110 73892
rect 59714 73836 59724 73892
rect 59780 73836 61404 73892
rect 61460 73836 61470 73892
rect 37986 73724 37996 73780
rect 38052 73724 40236 73780
rect 40292 73724 40302 73780
rect 41906 73724 41916 73780
rect 41972 73724 47068 73780
rect 47124 73724 47134 73780
rect 60050 73724 60060 73780
rect 60116 73724 60844 73780
rect 60900 73724 60910 73780
rect 19826 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20110 73724
rect 50546 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50830 73724
rect 32946 73612 32956 73668
rect 33012 73612 33740 73668
rect 33796 73612 34412 73668
rect 34468 73612 34478 73668
rect 38210 73612 38220 73668
rect 38276 73612 38668 73668
rect 38724 73612 38734 73668
rect 43250 73612 43260 73668
rect 43316 73612 47740 73668
rect 47796 73612 47806 73668
rect 55412 73556 55468 73668
rect 55524 73612 60732 73668
rect 60788 73612 60798 73668
rect 31602 73500 31612 73556
rect 31668 73500 32060 73556
rect 32116 73500 32126 73556
rect 32610 73500 32620 73556
rect 32676 73500 33628 73556
rect 33684 73500 33694 73556
rect 36642 73500 36652 73556
rect 36708 73500 40572 73556
rect 40628 73500 41468 73556
rect 41524 73500 41534 73556
rect 43474 73500 43484 73556
rect 43540 73500 43550 73556
rect 43810 73500 43820 73556
rect 43876 73500 45276 73556
rect 45332 73500 45342 73556
rect 45938 73500 45948 73556
rect 46004 73500 47068 73556
rect 47124 73500 47134 73556
rect 52434 73500 52444 73556
rect 52500 73500 53116 73556
rect 53172 73500 55468 73556
rect 56130 73500 56140 73556
rect 56196 73500 60508 73556
rect 60564 73500 60574 73556
rect 60946 73500 60956 73556
rect 61012 73500 61404 73556
rect 61460 73500 62300 73556
rect 62356 73500 62366 73556
rect 28466 73388 28476 73444
rect 28532 73388 30940 73444
rect 30996 73388 31276 73444
rect 31332 73388 31342 73444
rect 33394 73388 33404 73444
rect 33460 73388 34524 73444
rect 34580 73388 42364 73444
rect 42420 73388 42430 73444
rect 43484 73332 43540 73500
rect 60956 73444 61012 73500
rect 45378 73388 45388 73444
rect 45444 73388 45836 73444
rect 45892 73388 46508 73444
rect 46564 73388 46574 73444
rect 48738 73388 48748 73444
rect 48804 73388 50988 73444
rect 51044 73388 51772 73444
rect 51828 73388 51838 73444
rect 57810 73388 57820 73444
rect 57876 73388 58268 73444
rect 58324 73388 59500 73444
rect 59556 73388 59566 73444
rect 60274 73388 60284 73444
rect 60340 73388 61012 73444
rect 60284 73332 60340 73388
rect 37538 73276 37548 73332
rect 37604 73276 38220 73332
rect 38276 73276 38286 73332
rect 38658 73276 38668 73332
rect 38724 73276 40460 73332
rect 40516 73276 40526 73332
rect 43484 73276 45276 73332
rect 45332 73276 46396 73332
rect 46452 73276 49420 73332
rect 49476 73276 49486 73332
rect 52434 73276 52444 73332
rect 52500 73276 53564 73332
rect 53620 73276 57148 73332
rect 57204 73276 57214 73332
rect 58370 73276 58380 73332
rect 58436 73276 60340 73332
rect 43138 73164 43148 73220
rect 43204 73164 44268 73220
rect 44324 73164 45948 73220
rect 46004 73164 46014 73220
rect 48626 73164 48636 73220
rect 48692 73164 49644 73220
rect 49700 73164 49980 73220
rect 50036 73164 50046 73220
rect 42802 73052 42812 73108
rect 42868 73052 43596 73108
rect 43652 73052 43662 73108
rect 50082 73052 50092 73108
rect 50148 73052 50428 73108
rect 50484 73052 50988 73108
rect 51044 73052 51054 73108
rect 53890 73052 53900 73108
rect 53956 73052 54460 73108
rect 54516 73052 54908 73108
rect 54964 73052 55804 73108
rect 55860 73052 55870 73108
rect 41794 72940 41804 72996
rect 41860 72940 44604 72996
rect 44660 72940 44670 72996
rect 49858 72940 49868 72996
rect 49924 72940 52108 72996
rect 52164 72940 52174 72996
rect 56690 72940 56700 72996
rect 56756 72940 59388 72996
rect 59444 72940 59454 72996
rect 4466 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4750 72940
rect 35186 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35470 72940
rect 65906 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66190 72940
rect 30370 72716 30380 72772
rect 30436 72716 36540 72772
rect 36596 72716 36606 72772
rect 39106 72716 39116 72772
rect 39172 72716 40236 72772
rect 40292 72716 40302 72772
rect 55794 72716 55804 72772
rect 55860 72716 58828 72772
rect 58884 72716 58894 72772
rect 36194 72604 36204 72660
rect 36260 72604 42476 72660
rect 42532 72604 42542 72660
rect 54338 72604 54348 72660
rect 54404 72604 58604 72660
rect 58660 72604 58670 72660
rect 59042 72604 59052 72660
rect 59108 72604 60284 72660
rect 60340 72604 61964 72660
rect 62020 72604 62030 72660
rect 12898 72492 12908 72548
rect 12964 72492 35084 72548
rect 35140 72492 35150 72548
rect 41570 72492 41580 72548
rect 41636 72492 42588 72548
rect 42644 72492 44044 72548
rect 44100 72492 44110 72548
rect 44482 72492 44492 72548
rect 44548 72492 44940 72548
rect 44996 72492 45006 72548
rect 52098 72492 52108 72548
rect 52164 72492 52556 72548
rect 52612 72492 52780 72548
rect 52836 72492 53452 72548
rect 53508 72492 53518 72548
rect 55346 72492 55356 72548
rect 55412 72492 56028 72548
rect 56084 72492 56094 72548
rect 57026 72492 57036 72548
rect 57092 72492 59276 72548
rect 59332 72492 59342 72548
rect 44492 72436 44548 72492
rect 21410 72380 21420 72436
rect 21476 72380 34412 72436
rect 34468 72380 34478 72436
rect 35186 72380 35196 72436
rect 35252 72380 36204 72436
rect 36260 72380 36270 72436
rect 36530 72380 36540 72436
rect 36596 72380 37436 72436
rect 37492 72380 37502 72436
rect 37874 72380 37884 72436
rect 37940 72380 38892 72436
rect 38948 72380 41804 72436
rect 41860 72380 41870 72436
rect 43026 72380 43036 72436
rect 43092 72380 44548 72436
rect 48626 72380 48636 72436
rect 48692 72380 49420 72436
rect 49476 72380 49486 72436
rect 36418 72268 36428 72324
rect 36484 72268 36876 72324
rect 36932 72268 36942 72324
rect 41458 72268 41468 72324
rect 41524 72268 41534 72324
rect 41682 72268 41692 72324
rect 41748 72268 44156 72324
rect 44212 72268 45500 72324
rect 45556 72268 45566 72324
rect 48514 72268 48524 72324
rect 48580 72268 50876 72324
rect 50932 72268 51324 72324
rect 51380 72268 51884 72324
rect 51940 72268 51950 72324
rect 41468 72212 41524 72268
rect 37650 72156 37660 72212
rect 37716 72156 37996 72212
rect 38052 72156 38556 72212
rect 38612 72156 38780 72212
rect 38836 72156 38846 72212
rect 41234 72156 41244 72212
rect 41300 72156 41524 72212
rect 41906 72156 41916 72212
rect 41972 72156 45724 72212
rect 45780 72156 45790 72212
rect 45938 72156 45948 72212
rect 46004 72156 46172 72212
rect 46228 72156 46844 72212
rect 46900 72156 47292 72212
rect 47348 72156 47740 72212
rect 47796 72156 47806 72212
rect 55346 72156 55356 72212
rect 55412 72156 55916 72212
rect 55972 72156 55982 72212
rect 19826 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20110 72156
rect 41468 72100 41524 72156
rect 50546 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50830 72156
rect 36418 72044 36428 72100
rect 36484 72044 37548 72100
rect 37604 72044 37772 72100
rect 37828 72044 37838 72100
rect 41468 72044 43708 72100
rect 43764 72044 43774 72100
rect 45798 72044 45836 72100
rect 45892 72044 45902 72100
rect 37314 71932 37324 71988
rect 37380 71932 38332 71988
rect 38388 71932 42364 71988
rect 42420 71932 42430 71988
rect 43586 71932 43596 71988
rect 43652 71932 43820 71988
rect 43876 71932 43886 71988
rect 52882 71932 52892 71988
rect 52948 71932 53900 71988
rect 53956 71932 53966 71988
rect 34738 71820 34748 71876
rect 34804 71820 43708 71876
rect 43652 71764 43708 71820
rect 41234 71708 41244 71764
rect 41300 71708 42252 71764
rect 42308 71708 42924 71764
rect 42980 71708 42990 71764
rect 43652 71708 44604 71764
rect 44660 71708 44940 71764
rect 44996 71708 45006 71764
rect 50306 71708 50316 71764
rect 50372 71708 52556 71764
rect 52612 71708 52622 71764
rect 40114 71596 40124 71652
rect 40180 71596 41916 71652
rect 41972 71596 41982 71652
rect 56242 71484 56252 71540
rect 56308 71484 58268 71540
rect 58324 71484 58334 71540
rect 4466 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4750 71372
rect 35186 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35470 71372
rect 65906 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66190 71372
rect 36866 71260 36876 71316
rect 36932 71260 49532 71316
rect 49588 71260 49598 71316
rect 38770 71148 38780 71204
rect 38836 71148 39676 71204
rect 39732 71148 39742 71204
rect 34290 71036 34300 71092
rect 34356 71036 35308 71092
rect 35364 71036 36428 71092
rect 36484 71036 36494 71092
rect 40226 71036 40236 71092
rect 40292 71036 41020 71092
rect 41076 71036 42140 71092
rect 42196 71036 42206 71092
rect 43810 71036 43820 71092
rect 43876 71036 44492 71092
rect 44548 71036 44716 71092
rect 44772 71036 45388 71092
rect 45444 71036 45454 71092
rect 45938 71036 45948 71092
rect 46004 71036 49756 71092
rect 49812 71036 50876 71092
rect 50932 71036 50942 71092
rect 55412 71036 55692 71092
rect 55748 71036 56924 71092
rect 56980 71036 58940 71092
rect 58996 71036 59836 71092
rect 59892 71036 59902 71092
rect 38546 70924 38556 70980
rect 38612 70924 39676 70980
rect 39732 70924 39742 70980
rect 47842 70924 47852 70980
rect 47908 70924 48748 70980
rect 48804 70924 48814 70980
rect 55346 70924 55356 70980
rect 55412 70924 55468 71036
rect 38098 70812 38108 70868
rect 38164 70812 38780 70868
rect 38836 70812 40012 70868
rect 40068 70812 40460 70868
rect 40516 70812 40526 70868
rect 43362 70588 43372 70644
rect 43428 70588 43438 70644
rect 19826 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20110 70588
rect 43372 70532 43428 70588
rect 50546 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50830 70588
rect 31938 70476 31948 70532
rect 32004 70476 37380 70532
rect 43372 70476 45500 70532
rect 45556 70476 45566 70532
rect 46386 70476 46396 70532
rect 46452 70476 47852 70532
rect 47908 70476 47918 70532
rect 51314 70476 51324 70532
rect 51380 70476 52220 70532
rect 52276 70476 54124 70532
rect 54180 70476 60508 70532
rect 60564 70476 60574 70532
rect 37324 70420 37380 70476
rect 36306 70364 36316 70420
rect 36372 70364 37100 70420
rect 37156 70364 37166 70420
rect 37324 70364 48804 70420
rect 51762 70364 51772 70420
rect 51828 70364 52668 70420
rect 52724 70364 53564 70420
rect 53620 70364 53630 70420
rect 48748 70308 48804 70364
rect 37426 70252 37436 70308
rect 37492 70252 40348 70308
rect 40404 70252 40796 70308
rect 40852 70252 44828 70308
rect 44884 70252 46284 70308
rect 46340 70252 46350 70308
rect 48748 70252 53788 70308
rect 53844 70252 53854 70308
rect 37202 70140 37212 70196
rect 37268 70140 40236 70196
rect 40292 70140 40302 70196
rect 46162 70140 46172 70196
rect 46228 70140 47180 70196
rect 47236 70140 47246 70196
rect 4466 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4750 69804
rect 35186 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35470 69804
rect 65906 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66190 69804
rect 45154 69468 45164 69524
rect 45220 69468 46620 69524
rect 46676 69468 46686 69524
rect 50978 69468 50988 69524
rect 51044 69468 52780 69524
rect 52836 69468 52846 69524
rect 19826 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20110 69020
rect 50546 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50830 69020
rect 4466 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4750 68236
rect 35186 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35470 68236
rect 65906 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66190 68236
rect 19826 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20110 67452
rect 50546 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50830 67452
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 35186 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35470 66668
rect 65906 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66190 66668
rect 19826 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20110 65884
rect 50546 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50830 65884
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 35186 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35470 65100
rect 65906 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66190 65100
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 50546 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50830 64316
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 65906 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66190 63532
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 50546 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50830 62748
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 65906 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66190 61964
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 50546 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50830 61180
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 65906 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66190 60396
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 50546 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50830 59612
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 65906 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66190 58828
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 50546 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50830 58044
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 65906 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66190 57260
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 65906 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66190 55692
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 65906 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66190 54124
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 65906 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66190 52556
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 65906 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66190 50988
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 65906 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66190 49420
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 65906 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66190 47852
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 65906 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66190 46284
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 65906 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66190 44716
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 65906 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66190 43148
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 65906 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66190 41580
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 65906 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66190 40012
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 65906 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66190 38444
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 65906 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66190 36876
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 65906 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66190 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 65906 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66190 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 65906 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66190 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 65906 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66190 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 65906 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66190 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 65906 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66190 27468
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 65906 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66190 25900
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 65906 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66190 24332
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 65906 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66190 22764
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 65906 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66190 21196
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 65906 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66190 19628
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 65906 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66190 18060
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 65906 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66190 16492
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 65906 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66190 14924
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 65906 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66190 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 65906 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66190 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 65906 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66190 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 65906 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66190 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 65906 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66190 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 65906 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66190 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 73490 4396 73500 4452
rect 73556 4396 74060 4452
rect 74116 4396 74126 4452
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 65906 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66190 3948
rect 45042 3276 45052 3332
rect 45108 3276 45612 3332
rect 45668 3276 45678 3332
rect 47730 3276 47740 3332
rect 47796 3276 48860 3332
rect 48916 3276 48926 3332
rect 49746 3276 49756 3332
rect 49812 3276 50876 3332
rect 50932 3276 50942 3332
rect 51762 3276 51772 3332
rect 51828 3276 52780 3332
rect 52836 3276 52846 3332
rect 53106 3276 53116 3332
rect 53172 3276 54124 3332
rect 54180 3276 54190 3332
rect 54450 3276 54460 3332
rect 54516 3276 55468 3332
rect 55524 3276 55534 3332
rect 56466 3276 56476 3332
rect 56532 3276 57372 3332
rect 57428 3276 57438 3332
rect 58482 3276 58492 3332
rect 58548 3276 59388 3332
rect 59444 3276 59454 3332
rect 59826 3276 59836 3332
rect 59892 3276 60620 3332
rect 60676 3276 60686 3332
rect 61842 3276 61852 3332
rect 61908 3276 62636 3332
rect 62692 3276 62702 3332
rect 65314 3276 65324 3332
rect 65380 3276 65884 3332
rect 65940 3276 65950 3332
rect 66658 3276 66668 3332
rect 66724 3276 67228 3332
rect 67284 3276 67294 3332
rect 67890 3276 67900 3332
rect 67956 3276 69132 3332
rect 69188 3276 69198 3332
rect 71250 3276 71260 3332
rect 71316 3276 72380 3332
rect 72436 3276 72446 3332
rect 73266 3276 73276 3332
rect 73332 3276 74396 3332
rect 74452 3276 74462 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 69906 1820 69916 1876
rect 69972 1820 71148 1876
rect 71204 1820 71214 1876
rect 48402 1708 48412 1764
rect 48468 1708 49532 1764
rect 49588 1708 49598 1764
rect 68562 1708 68572 1764
rect 68628 1708 69804 1764
rect 69860 1708 69870 1764
rect 71922 1708 71932 1764
rect 71988 1708 73052 1764
rect 73108 1708 73118 1764
<< via3 >>
rect 19836 76804 19892 76860
rect 19940 76804 19996 76860
rect 20044 76804 20100 76860
rect 50556 76804 50612 76860
rect 50660 76804 50716 76860
rect 50764 76804 50820 76860
rect 4476 76020 4532 76076
rect 4580 76020 4636 76076
rect 4684 76020 4740 76076
rect 35196 76020 35252 76076
rect 35300 76020 35356 76076
rect 35404 76020 35460 76076
rect 65916 76020 65972 76076
rect 66020 76020 66076 76076
rect 66124 76020 66180 76076
rect 41692 75740 41748 75796
rect 19836 75236 19892 75292
rect 19940 75236 19996 75292
rect 20044 75236 20100 75292
rect 50556 75236 50612 75292
rect 50660 75236 50716 75292
rect 50764 75236 50820 75292
rect 51660 75180 51716 75236
rect 44604 75068 44660 75124
rect 41692 74844 41748 74900
rect 4476 74452 4532 74508
rect 4580 74452 4636 74508
rect 4684 74452 4740 74508
rect 35196 74452 35252 74508
rect 35300 74452 35356 74508
rect 35404 74452 35460 74508
rect 65916 74452 65972 74508
rect 66020 74452 66076 74508
rect 66124 74452 66180 74508
rect 51660 74284 51716 74340
rect 52220 74284 52276 74340
rect 45836 74060 45892 74116
rect 52220 73836 52276 73892
rect 19836 73668 19892 73724
rect 19940 73668 19996 73724
rect 20044 73668 20100 73724
rect 50556 73668 50612 73724
rect 50660 73668 50716 73724
rect 50764 73668 50820 73724
rect 4476 72884 4532 72940
rect 4580 72884 4636 72940
rect 4684 72884 4740 72940
rect 35196 72884 35252 72940
rect 35300 72884 35356 72940
rect 35404 72884 35460 72940
rect 65916 72884 65972 72940
rect 66020 72884 66076 72940
rect 66124 72884 66180 72940
rect 19836 72100 19892 72156
rect 19940 72100 19996 72156
rect 20044 72100 20100 72156
rect 50556 72100 50612 72156
rect 50660 72100 50716 72156
rect 50764 72100 50820 72156
rect 45836 72044 45892 72100
rect 44604 71708 44660 71764
rect 4476 71316 4532 71372
rect 4580 71316 4636 71372
rect 4684 71316 4740 71372
rect 35196 71316 35252 71372
rect 35300 71316 35356 71372
rect 35404 71316 35460 71372
rect 65916 71316 65972 71372
rect 66020 71316 66076 71372
rect 66124 71316 66180 71372
rect 19836 70532 19892 70588
rect 19940 70532 19996 70588
rect 20044 70532 20100 70588
rect 50556 70532 50612 70588
rect 50660 70532 50716 70588
rect 50764 70532 50820 70588
rect 4476 69748 4532 69804
rect 4580 69748 4636 69804
rect 4684 69748 4740 69804
rect 35196 69748 35252 69804
rect 35300 69748 35356 69804
rect 35404 69748 35460 69804
rect 65916 69748 65972 69804
rect 66020 69748 66076 69804
rect 66124 69748 66180 69804
rect 19836 68964 19892 69020
rect 19940 68964 19996 69020
rect 20044 68964 20100 69020
rect 50556 68964 50612 69020
rect 50660 68964 50716 69020
rect 50764 68964 50820 69020
rect 4476 68180 4532 68236
rect 4580 68180 4636 68236
rect 4684 68180 4740 68236
rect 35196 68180 35252 68236
rect 35300 68180 35356 68236
rect 35404 68180 35460 68236
rect 65916 68180 65972 68236
rect 66020 68180 66076 68236
rect 66124 68180 66180 68236
rect 19836 67396 19892 67452
rect 19940 67396 19996 67452
rect 20044 67396 20100 67452
rect 50556 67396 50612 67452
rect 50660 67396 50716 67452
rect 50764 67396 50820 67452
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 35196 66612 35252 66668
rect 35300 66612 35356 66668
rect 35404 66612 35460 66668
rect 65916 66612 65972 66668
rect 66020 66612 66076 66668
rect 66124 66612 66180 66668
rect 19836 65828 19892 65884
rect 19940 65828 19996 65884
rect 20044 65828 20100 65884
rect 50556 65828 50612 65884
rect 50660 65828 50716 65884
rect 50764 65828 50820 65884
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 35196 65044 35252 65100
rect 35300 65044 35356 65100
rect 35404 65044 35460 65100
rect 65916 65044 65972 65100
rect 66020 65044 66076 65100
rect 66124 65044 66180 65100
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 50556 64260 50612 64316
rect 50660 64260 50716 64316
rect 50764 64260 50820 64316
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 65916 63476 65972 63532
rect 66020 63476 66076 63532
rect 66124 63476 66180 63532
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 50556 62692 50612 62748
rect 50660 62692 50716 62748
rect 50764 62692 50820 62748
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 65916 61908 65972 61964
rect 66020 61908 66076 61964
rect 66124 61908 66180 61964
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 50556 61124 50612 61180
rect 50660 61124 50716 61180
rect 50764 61124 50820 61180
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 65916 60340 65972 60396
rect 66020 60340 66076 60396
rect 66124 60340 66180 60396
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 50556 59556 50612 59612
rect 50660 59556 50716 59612
rect 50764 59556 50820 59612
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 65916 58772 65972 58828
rect 66020 58772 66076 58828
rect 66124 58772 66180 58828
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 50556 57988 50612 58044
rect 50660 57988 50716 58044
rect 50764 57988 50820 58044
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 65916 57204 65972 57260
rect 66020 57204 66076 57260
rect 66124 57204 66180 57260
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 65916 55636 65972 55692
rect 66020 55636 66076 55692
rect 66124 55636 66180 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 65916 54068 65972 54124
rect 66020 54068 66076 54124
rect 66124 54068 66180 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 65916 52500 65972 52556
rect 66020 52500 66076 52556
rect 66124 52500 66180 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 65916 50932 65972 50988
rect 66020 50932 66076 50988
rect 66124 50932 66180 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 65916 49364 65972 49420
rect 66020 49364 66076 49420
rect 66124 49364 66180 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 65916 47796 65972 47852
rect 66020 47796 66076 47852
rect 66124 47796 66180 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 65916 46228 65972 46284
rect 66020 46228 66076 46284
rect 66124 46228 66180 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 65916 44660 65972 44716
rect 66020 44660 66076 44716
rect 66124 44660 66180 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 65916 43092 65972 43148
rect 66020 43092 66076 43148
rect 66124 43092 66180 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 65916 41524 65972 41580
rect 66020 41524 66076 41580
rect 66124 41524 66180 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 65916 39956 65972 40012
rect 66020 39956 66076 40012
rect 66124 39956 66180 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 65916 38388 65972 38444
rect 66020 38388 66076 38444
rect 66124 38388 66180 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 65916 36820 65972 36876
rect 66020 36820 66076 36876
rect 66124 36820 66180 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 65916 35252 65972 35308
rect 66020 35252 66076 35308
rect 66124 35252 66180 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 65916 33684 65972 33740
rect 66020 33684 66076 33740
rect 66124 33684 66180 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 65916 32116 65972 32172
rect 66020 32116 66076 32172
rect 66124 32116 66180 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 65916 30548 65972 30604
rect 66020 30548 66076 30604
rect 66124 30548 66180 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 65916 28980 65972 29036
rect 66020 28980 66076 29036
rect 66124 28980 66180 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 65916 27412 65972 27468
rect 66020 27412 66076 27468
rect 66124 27412 66180 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 65916 25844 65972 25900
rect 66020 25844 66076 25900
rect 66124 25844 66180 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 65916 24276 65972 24332
rect 66020 24276 66076 24332
rect 66124 24276 66180 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 65916 22708 65972 22764
rect 66020 22708 66076 22764
rect 66124 22708 66180 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 65916 21140 65972 21196
rect 66020 21140 66076 21196
rect 66124 21140 66180 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 65916 19572 65972 19628
rect 66020 19572 66076 19628
rect 66124 19572 66180 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 65916 18004 65972 18060
rect 66020 18004 66076 18060
rect 66124 18004 66180 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 65916 16436 65972 16492
rect 66020 16436 66076 16492
rect 66124 16436 66180 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 65916 14868 65972 14924
rect 66020 14868 66076 14924
rect 66124 14868 66180 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 65916 13300 65972 13356
rect 66020 13300 66076 13356
rect 66124 13300 66180 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 65916 11732 65972 11788
rect 66020 11732 66076 11788
rect 66124 11732 66180 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 65916 10164 65972 10220
rect 66020 10164 66076 10220
rect 66124 10164 66180 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 65916 8596 65972 8652
rect 66020 8596 66076 8652
rect 66124 8596 66180 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 65916 7028 65972 7084
rect 66020 7028 66076 7084
rect 66124 7028 66180 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 65916 5460 65972 5516
rect 66020 5460 66076 5516
rect 66124 5460 66180 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 65916 3892 65972 3948
rect 66020 3892 66076 3948
rect 66124 3892 66180 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 76076 4768 76892
rect 4448 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4768 76076
rect 4448 74508 4768 76020
rect 4448 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4768 74508
rect 4448 72940 4768 74452
rect 4448 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4768 72940
rect 4448 71372 4768 72884
rect 4448 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4768 71372
rect 4448 69804 4768 71316
rect 4448 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4768 69804
rect 4448 68236 4768 69748
rect 4448 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4768 68236
rect 4448 66668 4768 68180
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 76860 20128 76892
rect 19808 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20128 76860
rect 19808 75292 20128 76804
rect 19808 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20128 75292
rect 19808 73724 20128 75236
rect 19808 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20128 73724
rect 19808 72156 20128 73668
rect 19808 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20128 72156
rect 19808 70588 20128 72100
rect 19808 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20128 70588
rect 19808 69020 20128 70532
rect 19808 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20128 69020
rect 19808 67452 20128 68964
rect 19808 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20128 67452
rect 19808 65884 20128 67396
rect 19808 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20128 65884
rect 19808 64316 20128 65828
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 19808 61180 20128 62692
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19808 56476 20128 57988
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 76076 35488 76892
rect 35168 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35488 76076
rect 35168 74508 35488 76020
rect 50528 76860 50848 76892
rect 50528 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50848 76860
rect 41692 75796 41748 75806
rect 41692 74900 41748 75740
rect 50528 75292 50848 76804
rect 50528 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50848 75292
rect 65888 76076 66208 76892
rect 65888 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66208 76076
rect 41692 74834 41748 74844
rect 44604 75124 44660 75134
rect 35168 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35488 74508
rect 35168 72940 35488 74452
rect 35168 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35488 72940
rect 35168 71372 35488 72884
rect 44604 71764 44660 75068
rect 45836 74116 45892 74126
rect 45836 72100 45892 74060
rect 45836 72034 45892 72044
rect 50528 73724 50848 75236
rect 51660 75236 51716 75246
rect 51660 74340 51716 75180
rect 65888 74508 66208 76020
rect 65888 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66208 74508
rect 51660 74274 51716 74284
rect 52220 74340 52276 74350
rect 52220 73892 52276 74284
rect 52220 73826 52276 73836
rect 50528 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50848 73724
rect 50528 72156 50848 73668
rect 50528 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50848 72156
rect 44604 71698 44660 71708
rect 35168 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35488 71372
rect 35168 69804 35488 71316
rect 35168 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35488 69804
rect 35168 68236 35488 69748
rect 35168 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35488 68236
rect 35168 66668 35488 68180
rect 35168 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35488 66668
rect 35168 65100 35488 66612
rect 35168 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35488 65100
rect 35168 63532 35488 65044
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 35168 61964 35488 63476
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 35168 60396 35488 61908
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 35168 57260 35488 58772
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 70588 50848 72100
rect 50528 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50848 70588
rect 50528 69020 50848 70532
rect 50528 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50848 69020
rect 50528 67452 50848 68964
rect 50528 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50848 67452
rect 50528 65884 50848 67396
rect 50528 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50848 65884
rect 50528 64316 50848 65828
rect 50528 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50848 64316
rect 50528 62748 50848 64260
rect 50528 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50848 62748
rect 50528 61180 50848 62692
rect 50528 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50848 61180
rect 50528 59612 50848 61124
rect 50528 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50848 59612
rect 50528 58044 50848 59556
rect 50528 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50848 58044
rect 50528 56476 50848 57988
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 65888 72940 66208 74452
rect 65888 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66208 72940
rect 65888 71372 66208 72884
rect 65888 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66208 71372
rect 65888 69804 66208 71316
rect 65888 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66208 69804
rect 65888 68236 66208 69748
rect 65888 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66208 68236
rect 65888 66668 66208 68180
rect 65888 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66208 66668
rect 65888 65100 66208 66612
rect 65888 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66208 65100
rect 65888 63532 66208 65044
rect 65888 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66208 63532
rect 65888 61964 66208 63476
rect 65888 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66208 61964
rect 65888 60396 66208 61908
rect 65888 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66208 60396
rect 65888 58828 66208 60340
rect 65888 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66208 58828
rect 65888 57260 66208 58772
rect 65888 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66208 57260
rect 65888 55692 66208 57204
rect 65888 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66208 55692
rect 65888 54124 66208 55636
rect 65888 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66208 54124
rect 65888 52556 66208 54068
rect 65888 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66208 52556
rect 65888 50988 66208 52500
rect 65888 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66208 50988
rect 65888 49420 66208 50932
rect 65888 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66208 49420
rect 65888 47852 66208 49364
rect 65888 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66208 47852
rect 65888 46284 66208 47796
rect 65888 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66208 46284
rect 65888 44716 66208 46228
rect 65888 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66208 44716
rect 65888 43148 66208 44660
rect 65888 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66208 43148
rect 65888 41580 66208 43092
rect 65888 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66208 41580
rect 65888 40012 66208 41524
rect 65888 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66208 40012
rect 65888 38444 66208 39956
rect 65888 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66208 38444
rect 65888 36876 66208 38388
rect 65888 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66208 36876
rect 65888 35308 66208 36820
rect 65888 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66208 35308
rect 65888 33740 66208 35252
rect 65888 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66208 33740
rect 65888 32172 66208 33684
rect 65888 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66208 32172
rect 65888 30604 66208 32116
rect 65888 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66208 30604
rect 65888 29036 66208 30548
rect 65888 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66208 29036
rect 65888 27468 66208 28980
rect 65888 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66208 27468
rect 65888 25900 66208 27412
rect 65888 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66208 25900
rect 65888 24332 66208 25844
rect 65888 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66208 24332
rect 65888 22764 66208 24276
rect 65888 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66208 22764
rect 65888 21196 66208 22708
rect 65888 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66208 21196
rect 65888 19628 66208 21140
rect 65888 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66208 19628
rect 65888 18060 66208 19572
rect 65888 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66208 18060
rect 65888 16492 66208 18004
rect 65888 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66208 16492
rect 65888 14924 66208 16436
rect 65888 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66208 14924
rect 65888 13356 66208 14868
rect 65888 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66208 13356
rect 65888 11788 66208 13300
rect 65888 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66208 11788
rect 65888 10220 66208 11732
rect 65888 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66208 10220
rect 65888 8652 66208 10164
rect 65888 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66208 8652
rect 65888 7084 66208 8596
rect 65888 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66208 7084
rect 65888 5516 66208 7028
rect 65888 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66208 5516
rect 65888 3948 66208 5460
rect 65888 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66208 3948
rect 65888 3076 66208 3892
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__119__I dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 48720 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__123__A1
timestamp 1669390400
transform 1 0 47152 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__124__A1
timestamp 1669390400
transform -1 0 48272 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__124__A2
timestamp 1669390400
transform 1 0 46256 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__124__A3
timestamp 1669390400
transform 1 0 46704 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__125__A1
timestamp 1669390400
transform -1 0 47824 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__126__A1
timestamp 1669390400
transform 1 0 43792 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__I
timestamp 1669390400
transform 1 0 47376 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__A2
timestamp 1669390400
transform -1 0 46928 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__B2
timestamp 1669390400
transform 1 0 47824 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__129__A1
timestamp 1669390400
transform -1 0 48720 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__I
timestamp 1669390400
transform -1 0 37744 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__133__A2
timestamp 1669390400
transform -1 0 46480 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__134__A2
timestamp 1669390400
transform -1 0 40432 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__135__A2
timestamp 1669390400
transform -1 0 38192 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__136__I
timestamp 1669390400
transform 1 0 40768 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__138__A1
timestamp 1669390400
transform 1 0 41440 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__138__A3
timestamp 1669390400
transform 1 0 39760 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__141__A1
timestamp 1669390400
transform -1 0 44800 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__142__A1
timestamp 1669390400
transform -1 0 47376 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__147__I
timestamp 1669390400
transform 1 0 64512 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__150__A1
timestamp 1669390400
transform 1 0 62272 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__152__A1
timestamp 1669390400
transform 1 0 61936 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__152__A3
timestamp 1669390400
transform 1 0 59808 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__153__A1
timestamp 1669390400
transform 1 0 55440 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__154__A1
timestamp 1669390400
transform -1 0 52752 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__155__A1
timestamp 1669390400
transform 1 0 50848 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__156__I
timestamp 1669390400
transform 1 0 61376 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__157__A2
timestamp 1669390400
transform 1 0 61824 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__157__B2
timestamp 1669390400
transform 1 0 61264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__158__A1
timestamp 1669390400
transform 1 0 60256 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__159__A1
timestamp 1669390400
transform 1 0 55776 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__161__I
timestamp 1669390400
transform 1 0 55664 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__162__A2
timestamp 1669390400
transform 1 0 62832 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__167__A1
timestamp 1669390400
transform 1 0 58912 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__A1
timestamp 1669390400
transform 1 0 54656 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__170__A1
timestamp 1669390400
transform 1 0 54096 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__171__A1
timestamp 1669390400
transform -1 0 53648 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__171__B
timestamp 1669390400
transform -1 0 53200 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__176__I
timestamp 1669390400
transform 1 0 28784 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__A2
timestamp 1669390400
transform -1 0 50960 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__A2
timestamp 1669390400
transform -1 0 46032 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__B1
timestamp 1669390400
transform 1 0 52528 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__B2
timestamp 1669390400
transform 1 0 45024 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__I
timestamp 1669390400
transform -1 0 36176 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__I
timestamp 1669390400
transform 1 0 34720 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__A1
timestamp 1669390400
transform 1 0 37408 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__A1
timestamp 1669390400
transform 1 0 46256 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__I
timestamp 1669390400
transform -1 0 46256 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__A1
timestamp 1669390400
transform -1 0 33824 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__I
timestamp 1669390400
transform 1 0 62384 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__I
timestamp 1669390400
transform -1 0 29568 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__A2
timestamp 1669390400
transform -1 0 28224 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__A2
timestamp 1669390400
transform -1 0 28672 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__A1
timestamp 1669390400
transform -1 0 31024 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__A1
timestamp 1669390400
transform -1 0 29792 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__A2
timestamp 1669390400
transform -1 0 32032 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__A2
timestamp 1669390400
transform -1 0 39872 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__A2
timestamp 1669390400
transform 1 0 36400 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__I
timestamp 1669390400
transform -1 0 37744 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__I
timestamp 1669390400
transform -1 0 59696 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__S
timestamp 1669390400
transform 1 0 59024 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__A2
timestamp 1669390400
transform -1 0 33152 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__A1
timestamp 1669390400
transform -1 0 32704 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__A2
timestamp 1669390400
transform -1 0 34832 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__I
timestamp 1669390400
transform 1 0 38304 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__C
timestamp 1669390400
transform 1 0 49728 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__A2
timestamp 1669390400
transform -1 0 55104 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__C
timestamp 1669390400
transform -1 0 55552 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__A3
timestamp 1669390400
transform 1 0 55216 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__I
timestamp 1669390400
transform 1 0 33376 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__A1
timestamp 1669390400
transform 1 0 33824 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__A2
timestamp 1669390400
transform -1 0 36512 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__A1
timestamp 1669390400
transform -1 0 34048 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__A2
timestamp 1669390400
transform -1 0 35392 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__A1
timestamp 1669390400
transform 1 0 45360 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__A1
timestamp 1669390400
transform -1 0 40208 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__A1
timestamp 1669390400
transform -1 0 44352 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__B
timestamp 1669390400
transform 1 0 41216 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__A1
timestamp 1669390400
transform -1 0 52304 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__A1
timestamp 1669390400
transform 1 0 59696 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__A1
timestamp 1669390400
transform -1 0 51856 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__B
timestamp 1669390400
transform -1 0 51408 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__S
timestamp 1669390400
transform 1 0 49168 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__A1
timestamp 1669390400
transform -1 0 50512 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__A1
timestamp 1669390400
transform 1 0 50288 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__C
timestamp 1669390400
transform -1 0 49840 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__A2
timestamp 1669390400
transform -1 0 37184 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__B1
timestamp 1669390400
transform -1 0 36960 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__A2
timestamp 1669390400
transform 1 0 34272 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__I
timestamp 1669390400
transform -1 0 30016 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__A2
timestamp 1669390400
transform -1 0 33040 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1669390400
transform -1 0 1904 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform -1 0 38080 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1669390400
transform -1 0 40880 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1669390400
transform 1 0 45472 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1669390400
transform -1 0 46704 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1669390400
transform 1 0 48272 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1669390400
transform -1 0 48496 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1669390400
transform -1 0 52864 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1669390400
transform -1 0 52416 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1669390400
transform -1 0 54656 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1669390400
transform 1 0 63728 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1669390400
transform 1 0 64400 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1669390400
transform 1 0 63280 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1669390400
transform -1 0 62944 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1669390400
transform -1 0 65520 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1669390400
transform -1 0 68768 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1669390400
transform -1 0 69216 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1669390400
transform -1 0 70896 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1669390400
transform 1 0 73248 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1669390400
transform 1 0 77168 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1669390400
transform 1 0 78064 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output22_I
timestamp 1669390400
transform -1 0 7952 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output23_I
timestamp 1669390400
transform 1 0 24752 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output24_I
timestamp 1669390400
transform 1 0 26544 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output31_I
timestamp 1669390400
transform 1 0 12880 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output32_I
timestamp 1669390400
transform 1 0 15792 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output33_I
timestamp 1669390400
transform 1 0 17808 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output34_I
timestamp 1669390400
transform 1 0 19824 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output35_I
timestamp 1669390400
transform 1 0 20832 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output36_I
timestamp 1669390400
transform -1 0 24080 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_0_2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 3136
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_0_37 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5488 0 1 3136
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_0_45 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 6384 0 1 3136
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_0_53
timestamp 1669390400
transform 1 0 7280 0 1 3136
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 7728 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63
timestamp 1669390400
transform 1 0 8400 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1669390400
transform 1 0 9072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_0_72
timestamp 1669390400
transform 1 0 9408 0 1 3136
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80
timestamp 1669390400
transform 1 0 10304 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86
timestamp 1669390400
transform 1 0 10976 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92
timestamp 1669390400
transform 1 0 11648 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_98
timestamp 1669390400
transform 1 0 12320 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1669390400
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_0_107
timestamp 1669390400
transform 1 0 13328 0 1 3136
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_115
timestamp 1669390400
transform 1 0 14224 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_121
timestamp 1669390400
transform 1 0 14896 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_127
timestamp 1669390400
transform 1 0 15568 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_133
timestamp 1669390400
transform 1 0 16240 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1669390400
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_0_142
timestamp 1669390400
transform 1 0 17248 0 1 3136
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_150
timestamp 1669390400
transform 1 0 18144 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_156
timestamp 1669390400
transform 1 0 18816 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_162
timestamp 1669390400
transform 1 0 19488 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_168
timestamp 1669390400
transform 1 0 20160 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1669390400
transform 1 0 20832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_0_177
timestamp 1669390400
transform 1 0 21168 0 1 3136
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_185
timestamp 1669390400
transform 1 0 22064 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_191
timestamp 1669390400
transform 1 0 22736 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_197
timestamp 1669390400
transform 1 0 23408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_203
timestamp 1669390400
transform 1 0 24080 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1669390400
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_0_212
timestamp 1669390400
transform 1 0 25088 0 1 3136
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_220
timestamp 1669390400
transform 1 0 25984 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_226
timestamp 1669390400
transform 1 0 26656 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_232
timestamp 1669390400
transform 1 0 27328 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_238
timestamp 1669390400
transform 1 0 28000 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1669390400
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_0_247
timestamp 1669390400
transform 1 0 29008 0 1 3136
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_255
timestamp 1669390400
transform 1 0 29904 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_261
timestamp 1669390400
transform 1 0 30576 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_267
timestamp 1669390400
transform 1 0 31248 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_273
timestamp 1669390400
transform 1 0 31920 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1669390400
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_0_282
timestamp 1669390400
transform 1 0 32928 0 1 3136
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_290
timestamp 1669390400
transform 1 0 33824 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_296
timestamp 1669390400
transform 1 0 34496 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_302
timestamp 1669390400
transform 1 0 35168 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_308
timestamp 1669390400
transform 1 0 35840 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1669390400
transform 1 0 36512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_0_317
timestamp 1669390400
transform 1 0 36848 0 1 3136
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_325
timestamp 1669390400
transform 1 0 37744 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_331
timestamp 1669390400
transform 1 0 38416 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_337
timestamp 1669390400
transform 1 0 39088 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_343
timestamp 1669390400
transform 1 0 39760 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1669390400
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_352
timestamp 1669390400
transform 1 0 40768 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_354
timestamp 1669390400
transform 1 0 40992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_359
timestamp 1669390400
transform 1 0 41552 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_365
timestamp 1669390400
transform 1 0 42224 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_371
timestamp 1669390400
transform 1 0 42896 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_377
timestamp 1669390400
transform 1 0 43568 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_383
timestamp 1669390400
transform 1 0 44240 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_387
timestamp 1669390400
transform 1 0 44688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_392
timestamp 1669390400
transform 1 0 45248 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_398
timestamp 1669390400
transform 1 0 45920 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_404
timestamp 1669390400
transform 1 0 46592 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_410
timestamp 1669390400
transform 1 0 47264 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_0_416
timestamp 1669390400
transform 1 0 47936 0 1 3136
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_422
timestamp 1669390400
transform 1 0 48608 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_427
timestamp 1669390400
transform 1 0 49168 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_433
timestamp 1669390400
transform 1 0 49840 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_439
timestamp 1669390400
transform 1 0 50512 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_445
timestamp 1669390400
transform 1 0 51184 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_0_451
timestamp 1669390400
transform 1 0 51856 0 1 3136
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_457
timestamp 1669390400
transform 1 0 52528 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_462
timestamp 1669390400
transform 1 0 53088 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_468
timestamp 1669390400
transform 1 0 53760 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_474
timestamp 1669390400
transform 1 0 54432 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_480
timestamp 1669390400
transform 1 0 55104 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_0_486
timestamp 1669390400
transform 1 0 55776 0 1 3136
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_492
timestamp 1669390400
transform 1 0 56448 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_497
timestamp 1669390400
transform 1 0 57008 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_503
timestamp 1669390400
transform 1 0 57680 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_509
timestamp 1669390400
transform 1 0 58352 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_515
timestamp 1669390400
transform 1 0 59024 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_0_521
timestamp 1669390400
transform 1 0 59696 0 1 3136
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_527
timestamp 1669390400
transform 1 0 60368 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_532
timestamp 1669390400
transform 1 0 60928 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_538
timestamp 1669390400
transform 1 0 61600 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_544
timestamp 1669390400
transform 1 0 62272 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_550
timestamp 1669390400
transform 1 0 62944 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_0_556
timestamp 1669390400
transform 1 0 63616 0 1 3136
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_562
timestamp 1669390400
transform 1 0 64288 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_567
timestamp 1669390400
transform 1 0 64848 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_573
timestamp 1669390400
transform 1 0 65520 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_579
timestamp 1669390400
transform 1 0 66192 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_585
timestamp 1669390400
transform 1 0 66864 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_0_591
timestamp 1669390400
transform 1 0 67536 0 1 3136
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_597
timestamp 1669390400
transform 1 0 68208 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_602
timestamp 1669390400
transform 1 0 68768 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_608
timestamp 1669390400
transform 1 0 69440 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_614
timestamp 1669390400
transform 1 0 70112 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_620
timestamp 1669390400
transform 1 0 70784 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_0_626
timestamp 1669390400
transform 1 0 71456 0 1 3136
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_632
timestamp 1669390400
transform 1 0 72128 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_637
timestamp 1669390400
transform 1 0 72688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_643
timestamp 1669390400
transform 1 0 73360 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_649
timestamp 1669390400
transform 1 0 74032 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_0_655
timestamp 1669390400
transform 1 0 74704 0 1 3136
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_663
timestamp 1669390400
transform 1 0 75600 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_16  FILLER_0_667 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 76048 0 1 3136
box 0 -60 1792 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_0_683
timestamp 1669390400
transform 1 0 77840 0 1 3136
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_687
timestamp 1669390400
transform 1 0 78288 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_1_66
timestamp 1669390400
transform 1 0 8736 0 -1 4704
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1669390400
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_1_73
timestamp 1669390400
transform 1 0 9520 0 -1 4704
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_1_105
timestamp 1669390400
transform 1 0 13104 0 -1 4704
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_109
timestamp 1669390400
transform 1 0 13552 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_16  FILLER_1_115
timestamp 1669390400
transform 1 0 14224 0 -1 4704
box 0 -60 1792 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_1_131
timestamp 1669390400
transform 1 0 16016 0 -1 4704
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_139
timestamp 1669390400
transform 1 0 16912 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1669390400
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_144
timestamp 1669390400
transform 1 0 17472 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_146
timestamp 1669390400
transform 1 0 17696 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_1_151
timestamp 1669390400
transform 1 0 18256 0 -1 4704
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_16  FILLER_1_183
timestamp 1669390400
transform 1 0 21840 0 -1 4704
box 0 -60 1792 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_1_199
timestamp 1669390400
transform 1 0 23632 0 -1 4704
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_211
timestamp 1669390400
transform 1 0 24976 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_1_215
timestamp 1669390400
transform 1 0 25424 0 -1 4704
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_247
timestamp 1669390400
transform 1 0 29008 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_16  FILLER_1_253
timestamp 1669390400
transform 1 0 29680 0 -1 4704
box 0 -60 1792 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_1_269
timestamp 1669390400
transform 1 0 31472 0 -1 4704
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_281
timestamp 1669390400
transform 1 0 32816 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1669390400
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_1_286
timestamp 1669390400
transform 1 0 33376 0 -1 4704
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_318
timestamp 1669390400
transform 1 0 36960 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_1_323
timestamp 1669390400
transform 1 0 37520 0 -1 4704
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_357
timestamp 1669390400
transform 1 0 41328 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_1_421
timestamp 1669390400
transform 1 0 48496 0 -1 4704
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_425
timestamp 1669390400
transform 1 0 48944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_16  FILLER_1_428
timestamp 1669390400
transform 1 0 49280 0 -1 4704
box 0 -60 1792 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_444
timestamp 1669390400
transform 1 0 51072 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_1_449
timestamp 1669390400
transform 1 0 51632 0 -1 4704
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_1_485
timestamp 1669390400
transform 1 0 55664 0 -1 4704
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_1_493
timestamp 1669390400
transform 1 0 56560 0 -1 4704
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_16  FILLER_1_499
timestamp 1669390400
transform 1 0 57232 0 -1 4704
box 0 -60 1792 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_515
timestamp 1669390400
transform 1 0 59024 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_1_521
timestamp 1669390400
transform 1 0 59696 0 -1 4704
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_1_557
timestamp 1669390400
transform 1 0 63728 0 -1 4704
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_565
timestamp 1669390400
transform 1 0 64624 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_567
timestamp 1669390400
transform 1 0 64848 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_1_570
timestamp 1669390400
transform 1 0 65184 0 -1 4704
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_16  FILLER_1_602
timestamp 1669390400
transform 1 0 68768 0 -1 4704
box 0 -60 1792 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_618
timestamp 1669390400
transform 1 0 70560 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_16  FILLER_1_623
timestamp 1669390400
transform 1 0 71120 0 -1 4704
box 0 -60 1792 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_641
timestamp 1669390400
transform 1 0 73136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_646
timestamp 1669390400
transform 1 0 73696 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_1_652
timestamp 1669390400
transform 1 0 74368 0 -1 4704
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_1_684
timestamp 1669390400
transform 1 0 77952 0 -1 4704
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_2_2
timestamp 1669390400
transform 1 0 1568 0 1 4704
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1669390400
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1669390400
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_2_101
timestamp 1669390400
transform 1 0 12656 0 1 4704
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1669390400
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_108
timestamp 1669390400
transform 1 0 13440 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_2_172
timestamp 1669390400
transform 1 0 20608 0 1 4704
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1669390400
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_179
timestamp 1669390400
transform 1 0 21392 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_2_243
timestamp 1669390400
transform 1 0 28560 0 1 4704
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1669390400
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_250
timestamp 1669390400
transform 1 0 29344 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_2_314
timestamp 1669390400
transform 1 0 36512 0 1 4704
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1669390400
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_321
timestamp 1669390400
transform 1 0 37296 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_2_385
timestamp 1669390400
transform 1 0 44464 0 1 4704
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1669390400
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_392
timestamp 1669390400
transform 1 0 45248 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_2_456
timestamp 1669390400
transform 1 0 52416 0 1 4704
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_460
timestamp 1669390400
transform 1 0 52864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_463
timestamp 1669390400
transform 1 0 53200 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_2_527
timestamp 1669390400
transform 1 0 60368 0 1 4704
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_531
timestamp 1669390400
transform 1 0 60816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_534
timestamp 1669390400
transform 1 0 61152 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_2_598
timestamp 1669390400
transform 1 0 68320 0 1 4704
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_602
timestamp 1669390400
transform 1 0 68768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_605
timestamp 1669390400
transform 1 0 69104 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_2_669
timestamp 1669390400
transform 1 0 76272 0 1 4704
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_673
timestamp 1669390400
transform 1 0 76720 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_2_676
timestamp 1669390400
transform 1 0 77056 0 1 4704
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_2_684
timestamp 1669390400
transform 1 0 77952 0 1 4704
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1669390400
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_3_66
timestamp 1669390400
transform 1 0 8736 0 -1 6272
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1669390400
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_73
timestamp 1669390400
transform 1 0 9520 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_3_137
timestamp 1669390400
transform 1 0 16688 0 -1 6272
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1669390400
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_144
timestamp 1669390400
transform 1 0 17472 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_3_208
timestamp 1669390400
transform 1 0 24640 0 -1 6272
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1669390400
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_215
timestamp 1669390400
transform 1 0 25424 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_3_279
timestamp 1669390400
transform 1 0 32592 0 -1 6272
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1669390400
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_286
timestamp 1669390400
transform 1 0 33376 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_3_350
timestamp 1669390400
transform 1 0 40544 0 -1 6272
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1669390400
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_357
timestamp 1669390400
transform 1 0 41328 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_3_421
timestamp 1669390400
transform 1 0 48496 0 -1 6272
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_425
timestamp 1669390400
transform 1 0 48944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_428
timestamp 1669390400
transform 1 0 49280 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_3_492
timestamp 1669390400
transform 1 0 56448 0 -1 6272
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_496
timestamp 1669390400
transform 1 0 56896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_499
timestamp 1669390400
transform 1 0 57232 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_3_563
timestamp 1669390400
transform 1 0 64400 0 -1 6272
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_567
timestamp 1669390400
transform 1 0 64848 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_570
timestamp 1669390400
transform 1 0 65184 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_3_634
timestamp 1669390400
transform 1 0 72352 0 -1 6272
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_638
timestamp 1669390400
transform 1 0 72800 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_3_641
timestamp 1669390400
transform 1 0 73136 0 -1 6272
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_3_673
timestamp 1669390400
transform 1 0 76720 0 -1 6272
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_3_681
timestamp 1669390400
transform 1 0 77616 0 -1 6272
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_685
timestamp 1669390400
transform 1 0 78064 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_687
timestamp 1669390400
transform 1 0 78288 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_4_2
timestamp 1669390400
transform 1 0 1568 0 1 6272
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1669390400
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1669390400
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_4_101
timestamp 1669390400
transform 1 0 12656 0 1 6272
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1669390400
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_108
timestamp 1669390400
transform 1 0 13440 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_4_172
timestamp 1669390400
transform 1 0 20608 0 1 6272
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1669390400
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_179
timestamp 1669390400
transform 1 0 21392 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_4_243
timestamp 1669390400
transform 1 0 28560 0 1 6272
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1669390400
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_250
timestamp 1669390400
transform 1 0 29344 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_4_314
timestamp 1669390400
transform 1 0 36512 0 1 6272
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1669390400
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_321
timestamp 1669390400
transform 1 0 37296 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_4_385
timestamp 1669390400
transform 1 0 44464 0 1 6272
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1669390400
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_392
timestamp 1669390400
transform 1 0 45248 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_4_456
timestamp 1669390400
transform 1 0 52416 0 1 6272
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_460
timestamp 1669390400
transform 1 0 52864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_463
timestamp 1669390400
transform 1 0 53200 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_4_527
timestamp 1669390400
transform 1 0 60368 0 1 6272
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_531
timestamp 1669390400
transform 1 0 60816 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_534
timestamp 1669390400
transform 1 0 61152 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_4_598
timestamp 1669390400
transform 1 0 68320 0 1 6272
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_602
timestamp 1669390400
transform 1 0 68768 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_605
timestamp 1669390400
transform 1 0 69104 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_4_669
timestamp 1669390400
transform 1 0 76272 0 1 6272
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_673
timestamp 1669390400
transform 1 0 76720 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_4_676
timestamp 1669390400
transform 1 0 77056 0 1 6272
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_4_684
timestamp 1669390400
transform 1 0 77952 0 1 6272
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1669390400
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_5_66
timestamp 1669390400
transform 1 0 8736 0 -1 7840
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1669390400
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1669390400
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_5_137
timestamp 1669390400
transform 1 0 16688 0 -1 7840
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1669390400
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_144
timestamp 1669390400
transform 1 0 17472 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_5_208
timestamp 1669390400
transform 1 0 24640 0 -1 7840
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1669390400
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_215
timestamp 1669390400
transform 1 0 25424 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_5_279
timestamp 1669390400
transform 1 0 32592 0 -1 7840
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1669390400
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_286
timestamp 1669390400
transform 1 0 33376 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_5_350
timestamp 1669390400
transform 1 0 40544 0 -1 7840
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1669390400
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_357
timestamp 1669390400
transform 1 0 41328 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_5_421
timestamp 1669390400
transform 1 0 48496 0 -1 7840
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_425
timestamp 1669390400
transform 1 0 48944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_428
timestamp 1669390400
transform 1 0 49280 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_5_492
timestamp 1669390400
transform 1 0 56448 0 -1 7840
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1669390400
transform 1 0 56896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_499
timestamp 1669390400
transform 1 0 57232 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_5_563
timestamp 1669390400
transform 1 0 64400 0 -1 7840
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_567
timestamp 1669390400
transform 1 0 64848 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_570
timestamp 1669390400
transform 1 0 65184 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_5_634
timestamp 1669390400
transform 1 0 72352 0 -1 7840
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_638
timestamp 1669390400
transform 1 0 72800 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_5_641
timestamp 1669390400
transform 1 0 73136 0 -1 7840
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_5_673
timestamp 1669390400
transform 1 0 76720 0 -1 7840
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_5_681
timestamp 1669390400
transform 1 0 77616 0 -1 7840
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_685
timestamp 1669390400
transform 1 0 78064 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_687
timestamp 1669390400
transform 1 0 78288 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_6_2
timestamp 1669390400
transform 1 0 1568 0 1 7840
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1669390400
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1669390400
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_6_101
timestamp 1669390400
transform 1 0 12656 0 1 7840
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1669390400
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1669390400
transform 1 0 13440 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_6_172
timestamp 1669390400
transform 1 0 20608 0 1 7840
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1669390400
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_179
timestamp 1669390400
transform 1 0 21392 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_6_243
timestamp 1669390400
transform 1 0 28560 0 1 7840
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1669390400
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1669390400
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_6_314
timestamp 1669390400
transform 1 0 36512 0 1 7840
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1669390400
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1669390400
transform 1 0 37296 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_6_385
timestamp 1669390400
transform 1 0 44464 0 1 7840
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1669390400
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_392
timestamp 1669390400
transform 1 0 45248 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_6_456
timestamp 1669390400
transform 1 0 52416 0 1 7840
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_460
timestamp 1669390400
transform 1 0 52864 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_463
timestamp 1669390400
transform 1 0 53200 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_6_527
timestamp 1669390400
transform 1 0 60368 0 1 7840
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_531
timestamp 1669390400
transform 1 0 60816 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_534
timestamp 1669390400
transform 1 0 61152 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_6_598
timestamp 1669390400
transform 1 0 68320 0 1 7840
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_602
timestamp 1669390400
transform 1 0 68768 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_605
timestamp 1669390400
transform 1 0 69104 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_6_669
timestamp 1669390400
transform 1 0 76272 0 1 7840
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_673
timestamp 1669390400
transform 1 0 76720 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_6_676
timestamp 1669390400
transform 1 0 77056 0 1 7840
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_6_684
timestamp 1669390400
transform 1 0 77952 0 1 7840
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1669390400
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_7_66
timestamp 1669390400
transform 1 0 8736 0 -1 9408
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1669390400
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1669390400
transform 1 0 9520 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_7_137
timestamp 1669390400
transform 1 0 16688 0 -1 9408
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1669390400
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1669390400
transform 1 0 17472 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_7_208
timestamp 1669390400
transform 1 0 24640 0 -1 9408
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1669390400
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1669390400
transform 1 0 25424 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_7_279
timestamp 1669390400
transform 1 0 32592 0 -1 9408
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1669390400
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_286
timestamp 1669390400
transform 1 0 33376 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_7_350
timestamp 1669390400
transform 1 0 40544 0 -1 9408
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1669390400
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_357
timestamp 1669390400
transform 1 0 41328 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_7_421
timestamp 1669390400
transform 1 0 48496 0 -1 9408
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_425
timestamp 1669390400
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_428
timestamp 1669390400
transform 1 0 49280 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_7_492
timestamp 1669390400
transform 1 0 56448 0 -1 9408
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1669390400
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_499
timestamp 1669390400
transform 1 0 57232 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_7_563
timestamp 1669390400
transform 1 0 64400 0 -1 9408
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_567
timestamp 1669390400
transform 1 0 64848 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_570
timestamp 1669390400
transform 1 0 65184 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_7_634
timestamp 1669390400
transform 1 0 72352 0 -1 9408
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_638
timestamp 1669390400
transform 1 0 72800 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_7_641
timestamp 1669390400
transform 1 0 73136 0 -1 9408
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_7_673
timestamp 1669390400
transform 1 0 76720 0 -1 9408
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_7_681
timestamp 1669390400
transform 1 0 77616 0 -1 9408
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_685
timestamp 1669390400
transform 1 0 78064 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_687
timestamp 1669390400
transform 1 0 78288 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_8_2
timestamp 1669390400
transform 1 0 1568 0 1 9408
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1669390400
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1669390400
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_8_101
timestamp 1669390400
transform 1 0 12656 0 1 9408
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1669390400
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1669390400
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_8_172
timestamp 1669390400
transform 1 0 20608 0 1 9408
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1669390400
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1669390400
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_8_243
timestamp 1669390400
transform 1 0 28560 0 1 9408
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1669390400
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1669390400
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_8_314
timestamp 1669390400
transform 1 0 36512 0 1 9408
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1669390400
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_321
timestamp 1669390400
transform 1 0 37296 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_8_385
timestamp 1669390400
transform 1 0 44464 0 1 9408
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1669390400
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_392
timestamp 1669390400
transform 1 0 45248 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_8_456
timestamp 1669390400
transform 1 0 52416 0 1 9408
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1669390400
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_463
timestamp 1669390400
transform 1 0 53200 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_8_527
timestamp 1669390400
transform 1 0 60368 0 1 9408
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_531
timestamp 1669390400
transform 1 0 60816 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_534
timestamp 1669390400
transform 1 0 61152 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_8_598
timestamp 1669390400
transform 1 0 68320 0 1 9408
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_602
timestamp 1669390400
transform 1 0 68768 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_605
timestamp 1669390400
transform 1 0 69104 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_8_669
timestamp 1669390400
transform 1 0 76272 0 1 9408
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_673
timestamp 1669390400
transform 1 0 76720 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_8_676
timestamp 1669390400
transform 1 0 77056 0 1 9408
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_8_684
timestamp 1669390400
transform 1 0 77952 0 1 9408
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1669390400
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_9_66
timestamp 1669390400
transform 1 0 8736 0 -1 10976
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1669390400
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1669390400
transform 1 0 9520 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_9_137
timestamp 1669390400
transform 1 0 16688 0 -1 10976
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1669390400
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1669390400
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_9_208
timestamp 1669390400
transform 1 0 24640 0 -1 10976
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1669390400
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1669390400
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_9_279
timestamp 1669390400
transform 1 0 32592 0 -1 10976
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1669390400
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_286
timestamp 1669390400
transform 1 0 33376 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_9_350
timestamp 1669390400
transform 1 0 40544 0 -1 10976
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1669390400
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_357
timestamp 1669390400
transform 1 0 41328 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_9_421
timestamp 1669390400
transform 1 0 48496 0 -1 10976
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_425
timestamp 1669390400
transform 1 0 48944 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_428
timestamp 1669390400
transform 1 0 49280 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_9_492
timestamp 1669390400
transform 1 0 56448 0 -1 10976
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1669390400
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_499
timestamp 1669390400
transform 1 0 57232 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_9_563
timestamp 1669390400
transform 1 0 64400 0 -1 10976
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_567
timestamp 1669390400
transform 1 0 64848 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_570
timestamp 1669390400
transform 1 0 65184 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_9_634
timestamp 1669390400
transform 1 0 72352 0 -1 10976
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_638
timestamp 1669390400
transform 1 0 72800 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_9_641
timestamp 1669390400
transform 1 0 73136 0 -1 10976
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_9_673
timestamp 1669390400
transform 1 0 76720 0 -1 10976
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_9_681
timestamp 1669390400
transform 1 0 77616 0 -1 10976
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_685
timestamp 1669390400
transform 1 0 78064 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_687
timestamp 1669390400
transform 1 0 78288 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_10_2
timestamp 1669390400
transform 1 0 1568 0 1 10976
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1669390400
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1669390400
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_10_101
timestamp 1669390400
transform 1 0 12656 0 1 10976
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1669390400
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1669390400
transform 1 0 13440 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_10_172
timestamp 1669390400
transform 1 0 20608 0 1 10976
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1669390400
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1669390400
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_10_243
timestamp 1669390400
transform 1 0 28560 0 1 10976
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1669390400
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1669390400
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_10_314
timestamp 1669390400
transform 1 0 36512 0 1 10976
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1669390400
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_321
timestamp 1669390400
transform 1 0 37296 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_10_385
timestamp 1669390400
transform 1 0 44464 0 1 10976
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1669390400
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_392
timestamp 1669390400
transform 1 0 45248 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_10_456
timestamp 1669390400
transform 1 0 52416 0 1 10976
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_460
timestamp 1669390400
transform 1 0 52864 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_463
timestamp 1669390400
transform 1 0 53200 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_10_527
timestamp 1669390400
transform 1 0 60368 0 1 10976
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_531
timestamp 1669390400
transform 1 0 60816 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_534
timestamp 1669390400
transform 1 0 61152 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_10_598
timestamp 1669390400
transform 1 0 68320 0 1 10976
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_602
timestamp 1669390400
transform 1 0 68768 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_605
timestamp 1669390400
transform 1 0 69104 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_10_669
timestamp 1669390400
transform 1 0 76272 0 1 10976
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_673
timestamp 1669390400
transform 1 0 76720 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_10_676
timestamp 1669390400
transform 1 0 77056 0 1 10976
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_10_684
timestamp 1669390400
transform 1 0 77952 0 1 10976
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1669390400
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_11_66
timestamp 1669390400
transform 1 0 8736 0 -1 12544
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1669390400
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1669390400
transform 1 0 9520 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_11_137
timestamp 1669390400
transform 1 0 16688 0 -1 12544
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1669390400
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1669390400
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_11_208
timestamp 1669390400
transform 1 0 24640 0 -1 12544
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1669390400
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1669390400
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_11_279
timestamp 1669390400
transform 1 0 32592 0 -1 12544
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1669390400
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_286
timestamp 1669390400
transform 1 0 33376 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_11_350
timestamp 1669390400
transform 1 0 40544 0 -1 12544
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1669390400
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_357
timestamp 1669390400
transform 1 0 41328 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_11_421
timestamp 1669390400
transform 1 0 48496 0 -1 12544
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_425
timestamp 1669390400
transform 1 0 48944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_428
timestamp 1669390400
transform 1 0 49280 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_11_492
timestamp 1669390400
transform 1 0 56448 0 -1 12544
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_496
timestamp 1669390400
transform 1 0 56896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_499
timestamp 1669390400
transform 1 0 57232 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_11_563
timestamp 1669390400
transform 1 0 64400 0 -1 12544
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_567
timestamp 1669390400
transform 1 0 64848 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_570
timestamp 1669390400
transform 1 0 65184 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_11_634
timestamp 1669390400
transform 1 0 72352 0 -1 12544
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_638
timestamp 1669390400
transform 1 0 72800 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_11_641
timestamp 1669390400
transform 1 0 73136 0 -1 12544
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_11_673
timestamp 1669390400
transform 1 0 76720 0 -1 12544
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_11_681
timestamp 1669390400
transform 1 0 77616 0 -1 12544
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_685
timestamp 1669390400
transform 1 0 78064 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_687
timestamp 1669390400
transform 1 0 78288 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_12_2
timestamp 1669390400
transform 1 0 1568 0 1 12544
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1669390400
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1669390400
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_12_101
timestamp 1669390400
transform 1 0 12656 0 1 12544
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1669390400
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1669390400
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_12_172
timestamp 1669390400
transform 1 0 20608 0 1 12544
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1669390400
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1669390400
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_12_243
timestamp 1669390400
transform 1 0 28560 0 1 12544
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1669390400
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1669390400
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_12_314
timestamp 1669390400
transform 1 0 36512 0 1 12544
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1669390400
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1669390400
transform 1 0 37296 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_12_385
timestamp 1669390400
transform 1 0 44464 0 1 12544
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1669390400
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_392
timestamp 1669390400
transform 1 0 45248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_12_456
timestamp 1669390400
transform 1 0 52416 0 1 12544
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1669390400
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_463
timestamp 1669390400
transform 1 0 53200 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_12_527
timestamp 1669390400
transform 1 0 60368 0 1 12544
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_531
timestamp 1669390400
transform 1 0 60816 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_534
timestamp 1669390400
transform 1 0 61152 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_12_598
timestamp 1669390400
transform 1 0 68320 0 1 12544
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_602
timestamp 1669390400
transform 1 0 68768 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_605
timestamp 1669390400
transform 1 0 69104 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_12_669
timestamp 1669390400
transform 1 0 76272 0 1 12544
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_673
timestamp 1669390400
transform 1 0 76720 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_12_676
timestamp 1669390400
transform 1 0 77056 0 1 12544
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_12_684
timestamp 1669390400
transform 1 0 77952 0 1 12544
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1669390400
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_13_66
timestamp 1669390400
transform 1 0 8736 0 -1 14112
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1669390400
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_73
timestamp 1669390400
transform 1 0 9520 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_13_137
timestamp 1669390400
transform 1 0 16688 0 -1 14112
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1669390400
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1669390400
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_13_208
timestamp 1669390400
transform 1 0 24640 0 -1 14112
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1669390400
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1669390400
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_13_279
timestamp 1669390400
transform 1 0 32592 0 -1 14112
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1669390400
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1669390400
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_13_350
timestamp 1669390400
transform 1 0 40544 0 -1 14112
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1669390400
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_357
timestamp 1669390400
transform 1 0 41328 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_13_421
timestamp 1669390400
transform 1 0 48496 0 -1 14112
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_425
timestamp 1669390400
transform 1 0 48944 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_428
timestamp 1669390400
transform 1 0 49280 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_13_492
timestamp 1669390400
transform 1 0 56448 0 -1 14112
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_496
timestamp 1669390400
transform 1 0 56896 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_499
timestamp 1669390400
transform 1 0 57232 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_13_563
timestamp 1669390400
transform 1 0 64400 0 -1 14112
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_567
timestamp 1669390400
transform 1 0 64848 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_570
timestamp 1669390400
transform 1 0 65184 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_13_634
timestamp 1669390400
transform 1 0 72352 0 -1 14112
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_638
timestamp 1669390400
transform 1 0 72800 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_13_641
timestamp 1669390400
transform 1 0 73136 0 -1 14112
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_13_673
timestamp 1669390400
transform 1 0 76720 0 -1 14112
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_13_681
timestamp 1669390400
transform 1 0 77616 0 -1 14112
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_685
timestamp 1669390400
transform 1 0 78064 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_687
timestamp 1669390400
transform 1 0 78288 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_14_2
timestamp 1669390400
transform 1 0 1568 0 1 14112
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1669390400
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1669390400
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_14_101
timestamp 1669390400
transform 1 0 12656 0 1 14112
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1669390400
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1669390400
transform 1 0 13440 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_14_172
timestamp 1669390400
transform 1 0 20608 0 1 14112
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1669390400
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1669390400
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_14_243
timestamp 1669390400
transform 1 0 28560 0 1 14112
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1669390400
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1669390400
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_14_314
timestamp 1669390400
transform 1 0 36512 0 1 14112
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1669390400
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1669390400
transform 1 0 37296 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_14_385
timestamp 1669390400
transform 1 0 44464 0 1 14112
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1669390400
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_392
timestamp 1669390400
transform 1 0 45248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_14_456
timestamp 1669390400
transform 1 0 52416 0 1 14112
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_460
timestamp 1669390400
transform 1 0 52864 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_463
timestamp 1669390400
transform 1 0 53200 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_14_527
timestamp 1669390400
transform 1 0 60368 0 1 14112
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_531
timestamp 1669390400
transform 1 0 60816 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_534
timestamp 1669390400
transform 1 0 61152 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_14_598
timestamp 1669390400
transform 1 0 68320 0 1 14112
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_602
timestamp 1669390400
transform 1 0 68768 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_605
timestamp 1669390400
transform 1 0 69104 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_14_669
timestamp 1669390400
transform 1 0 76272 0 1 14112
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_673
timestamp 1669390400
transform 1 0 76720 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_14_676
timestamp 1669390400
transform 1 0 77056 0 1 14112
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_14_684
timestamp 1669390400
transform 1 0 77952 0 1 14112
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1669390400
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_15_66
timestamp 1669390400
transform 1 0 8736 0 -1 15680
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1669390400
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1669390400
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_15_137
timestamp 1669390400
transform 1 0 16688 0 -1 15680
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1669390400
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1669390400
transform 1 0 17472 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_15_208
timestamp 1669390400
transform 1 0 24640 0 -1 15680
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1669390400
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1669390400
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_15_279
timestamp 1669390400
transform 1 0 32592 0 -1 15680
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1669390400
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1669390400
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_15_350
timestamp 1669390400
transform 1 0 40544 0 -1 15680
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1669390400
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_357
timestamp 1669390400
transform 1 0 41328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_15_421
timestamp 1669390400
transform 1 0 48496 0 -1 15680
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1669390400
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_428
timestamp 1669390400
transform 1 0 49280 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_15_492
timestamp 1669390400
transform 1 0 56448 0 -1 15680
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_496
timestamp 1669390400
transform 1 0 56896 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_499
timestamp 1669390400
transform 1 0 57232 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_15_563
timestamp 1669390400
transform 1 0 64400 0 -1 15680
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_567
timestamp 1669390400
transform 1 0 64848 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_570
timestamp 1669390400
transform 1 0 65184 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_15_634
timestamp 1669390400
transform 1 0 72352 0 -1 15680
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_638
timestamp 1669390400
transform 1 0 72800 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_15_641
timestamp 1669390400
transform 1 0 73136 0 -1 15680
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_15_673
timestamp 1669390400
transform 1 0 76720 0 -1 15680
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_15_681
timestamp 1669390400
transform 1 0 77616 0 -1 15680
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_685
timestamp 1669390400
transform 1 0 78064 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_687
timestamp 1669390400
transform 1 0 78288 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_16_2
timestamp 1669390400
transform 1 0 1568 0 1 15680
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1669390400
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1669390400
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_16_101
timestamp 1669390400
transform 1 0 12656 0 1 15680
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1669390400
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_108
timestamp 1669390400
transform 1 0 13440 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_16_172
timestamp 1669390400
transform 1 0 20608 0 1 15680
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1669390400
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_179
timestamp 1669390400
transform 1 0 21392 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_16_243
timestamp 1669390400
transform 1 0 28560 0 1 15680
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1669390400
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1669390400
transform 1 0 29344 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_16_314
timestamp 1669390400
transform 1 0 36512 0 1 15680
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1669390400
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_321
timestamp 1669390400
transform 1 0 37296 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_16_385
timestamp 1669390400
transform 1 0 44464 0 1 15680
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1669390400
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_392
timestamp 1669390400
transform 1 0 45248 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_16_456
timestamp 1669390400
transform 1 0 52416 0 1 15680
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_460
timestamp 1669390400
transform 1 0 52864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_463
timestamp 1669390400
transform 1 0 53200 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_16_527
timestamp 1669390400
transform 1 0 60368 0 1 15680
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_531
timestamp 1669390400
transform 1 0 60816 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_534
timestamp 1669390400
transform 1 0 61152 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_16_598
timestamp 1669390400
transform 1 0 68320 0 1 15680
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_602
timestamp 1669390400
transform 1 0 68768 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_605
timestamp 1669390400
transform 1 0 69104 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_16_669
timestamp 1669390400
transform 1 0 76272 0 1 15680
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_673
timestamp 1669390400
transform 1 0 76720 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_16_676
timestamp 1669390400
transform 1 0 77056 0 1 15680
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_16_684
timestamp 1669390400
transform 1 0 77952 0 1 15680
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_2
timestamp 1669390400
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_17_66
timestamp 1669390400
transform 1 0 8736 0 -1 17248
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1669390400
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_73
timestamp 1669390400
transform 1 0 9520 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_17_137
timestamp 1669390400
transform 1 0 16688 0 -1 17248
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1669390400
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_144
timestamp 1669390400
transform 1 0 17472 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_17_208
timestamp 1669390400
transform 1 0 24640 0 -1 17248
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1669390400
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_215
timestamp 1669390400
transform 1 0 25424 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_17_279
timestamp 1669390400
transform 1 0 32592 0 -1 17248
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1669390400
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_286
timestamp 1669390400
transform 1 0 33376 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_17_350
timestamp 1669390400
transform 1 0 40544 0 -1 17248
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1669390400
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_357
timestamp 1669390400
transform 1 0 41328 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_17_421
timestamp 1669390400
transform 1 0 48496 0 -1 17248
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_425
timestamp 1669390400
transform 1 0 48944 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_428
timestamp 1669390400
transform 1 0 49280 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_17_492
timestamp 1669390400
transform 1 0 56448 0 -1 17248
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_496
timestamp 1669390400
transform 1 0 56896 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_499
timestamp 1669390400
transform 1 0 57232 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_17_563
timestamp 1669390400
transform 1 0 64400 0 -1 17248
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_567
timestamp 1669390400
transform 1 0 64848 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_570
timestamp 1669390400
transform 1 0 65184 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_17_634
timestamp 1669390400
transform 1 0 72352 0 -1 17248
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_638
timestamp 1669390400
transform 1 0 72800 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_17_641
timestamp 1669390400
transform 1 0 73136 0 -1 17248
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_17_673
timestamp 1669390400
transform 1 0 76720 0 -1 17248
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_17_681
timestamp 1669390400
transform 1 0 77616 0 -1 17248
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_685
timestamp 1669390400
transform 1 0 78064 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_687
timestamp 1669390400
transform 1 0 78288 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_18_2
timestamp 1669390400
transform 1 0 1568 0 1 17248
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1669390400
transform 1 0 5152 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1669390400
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_18_101
timestamp 1669390400
transform 1 0 12656 0 1 17248
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1669390400
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_108
timestamp 1669390400
transform 1 0 13440 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_18_172
timestamp 1669390400
transform 1 0 20608 0 1 17248
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1669390400
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_179
timestamp 1669390400
transform 1 0 21392 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_18_243
timestamp 1669390400
transform 1 0 28560 0 1 17248
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1669390400
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1669390400
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_18_314
timestamp 1669390400
transform 1 0 36512 0 1 17248
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1669390400
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_321
timestamp 1669390400
transform 1 0 37296 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_18_385
timestamp 1669390400
transform 1 0 44464 0 1 17248
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1669390400
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_392
timestamp 1669390400
transform 1 0 45248 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_18_456
timestamp 1669390400
transform 1 0 52416 0 1 17248
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_460
timestamp 1669390400
transform 1 0 52864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_463
timestamp 1669390400
transform 1 0 53200 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_18_527
timestamp 1669390400
transform 1 0 60368 0 1 17248
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_531
timestamp 1669390400
transform 1 0 60816 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_534
timestamp 1669390400
transform 1 0 61152 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_18_598
timestamp 1669390400
transform 1 0 68320 0 1 17248
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_602
timestamp 1669390400
transform 1 0 68768 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_605
timestamp 1669390400
transform 1 0 69104 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_18_669
timestamp 1669390400
transform 1 0 76272 0 1 17248
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_673
timestamp 1669390400
transform 1 0 76720 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_18_676
timestamp 1669390400
transform 1 0 77056 0 1 17248
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_18_684
timestamp 1669390400
transform 1 0 77952 0 1 17248
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_2
timestamp 1669390400
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_19_66
timestamp 1669390400
transform 1 0 8736 0 -1 18816
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1669390400
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1669390400
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_19_137
timestamp 1669390400
transform 1 0 16688 0 -1 18816
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1669390400
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_144
timestamp 1669390400
transform 1 0 17472 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_19_208
timestamp 1669390400
transform 1 0 24640 0 -1 18816
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1669390400
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1669390400
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_19_279
timestamp 1669390400
transform 1 0 32592 0 -1 18816
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1669390400
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1669390400
transform 1 0 33376 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_19_350
timestamp 1669390400
transform 1 0 40544 0 -1 18816
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1669390400
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_357
timestamp 1669390400
transform 1 0 41328 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_19_421
timestamp 1669390400
transform 1 0 48496 0 -1 18816
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_425
timestamp 1669390400
transform 1 0 48944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_428
timestamp 1669390400
transform 1 0 49280 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_19_492
timestamp 1669390400
transform 1 0 56448 0 -1 18816
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_496
timestamp 1669390400
transform 1 0 56896 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_499
timestamp 1669390400
transform 1 0 57232 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_19_563
timestamp 1669390400
transform 1 0 64400 0 -1 18816
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_567
timestamp 1669390400
transform 1 0 64848 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_570
timestamp 1669390400
transform 1 0 65184 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_19_634
timestamp 1669390400
transform 1 0 72352 0 -1 18816
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_638
timestamp 1669390400
transform 1 0 72800 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_19_641
timestamp 1669390400
transform 1 0 73136 0 -1 18816
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_19_673
timestamp 1669390400
transform 1 0 76720 0 -1 18816
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_19_681
timestamp 1669390400
transform 1 0 77616 0 -1 18816
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_685
timestamp 1669390400
transform 1 0 78064 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_687
timestamp 1669390400
transform 1 0 78288 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_20_2
timestamp 1669390400
transform 1 0 1568 0 1 18816
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1669390400
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1669390400
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_20_101
timestamp 1669390400
transform 1 0 12656 0 1 18816
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1669390400
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1669390400
transform 1 0 13440 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_20_172
timestamp 1669390400
transform 1 0 20608 0 1 18816
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1669390400
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_179
timestamp 1669390400
transform 1 0 21392 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_20_243
timestamp 1669390400
transform 1 0 28560 0 1 18816
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1669390400
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1669390400
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_20_314
timestamp 1669390400
transform 1 0 36512 0 1 18816
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1669390400
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_321
timestamp 1669390400
transform 1 0 37296 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_20_385
timestamp 1669390400
transform 1 0 44464 0 1 18816
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1669390400
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_392
timestamp 1669390400
transform 1 0 45248 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_20_456
timestamp 1669390400
transform 1 0 52416 0 1 18816
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_460
timestamp 1669390400
transform 1 0 52864 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_463
timestamp 1669390400
transform 1 0 53200 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_20_527
timestamp 1669390400
transform 1 0 60368 0 1 18816
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_531
timestamp 1669390400
transform 1 0 60816 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_534
timestamp 1669390400
transform 1 0 61152 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_20_598
timestamp 1669390400
transform 1 0 68320 0 1 18816
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_602
timestamp 1669390400
transform 1 0 68768 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_605
timestamp 1669390400
transform 1 0 69104 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_20_669
timestamp 1669390400
transform 1 0 76272 0 1 18816
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_673
timestamp 1669390400
transform 1 0 76720 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_20_676
timestamp 1669390400
transform 1 0 77056 0 1 18816
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_20_684
timestamp 1669390400
transform 1 0 77952 0 1 18816
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1669390400
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_21_66
timestamp 1669390400
transform 1 0 8736 0 -1 20384
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1669390400
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1669390400
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_21_137
timestamp 1669390400
transform 1 0 16688 0 -1 20384
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1669390400
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_144
timestamp 1669390400
transform 1 0 17472 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_21_208
timestamp 1669390400
transform 1 0 24640 0 -1 20384
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1669390400
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1669390400
transform 1 0 25424 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_21_279
timestamp 1669390400
transform 1 0 32592 0 -1 20384
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1669390400
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1669390400
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_21_350
timestamp 1669390400
transform 1 0 40544 0 -1 20384
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1669390400
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_357
timestamp 1669390400
transform 1 0 41328 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_21_421
timestamp 1669390400
transform 1 0 48496 0 -1 20384
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_425
timestamp 1669390400
transform 1 0 48944 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_428
timestamp 1669390400
transform 1 0 49280 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_21_492
timestamp 1669390400
transform 1 0 56448 0 -1 20384
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_496
timestamp 1669390400
transform 1 0 56896 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_499
timestamp 1669390400
transform 1 0 57232 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_21_563
timestamp 1669390400
transform 1 0 64400 0 -1 20384
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_567
timestamp 1669390400
transform 1 0 64848 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_570
timestamp 1669390400
transform 1 0 65184 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_21_634
timestamp 1669390400
transform 1 0 72352 0 -1 20384
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_638
timestamp 1669390400
transform 1 0 72800 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_21_641
timestamp 1669390400
transform 1 0 73136 0 -1 20384
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_21_673
timestamp 1669390400
transform 1 0 76720 0 -1 20384
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_21_681
timestamp 1669390400
transform 1 0 77616 0 -1 20384
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_685
timestamp 1669390400
transform 1 0 78064 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_687
timestamp 1669390400
transform 1 0 78288 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_22_2
timestamp 1669390400
transform 1 0 1568 0 1 20384
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1669390400
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1669390400
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_22_101
timestamp 1669390400
transform 1 0 12656 0 1 20384
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1669390400
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1669390400
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_22_172
timestamp 1669390400
transform 1 0 20608 0 1 20384
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1669390400
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1669390400
transform 1 0 21392 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_22_243
timestamp 1669390400
transform 1 0 28560 0 1 20384
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1669390400
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1669390400
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_22_314
timestamp 1669390400
transform 1 0 36512 0 1 20384
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1669390400
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_321
timestamp 1669390400
transform 1 0 37296 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_22_385
timestamp 1669390400
transform 1 0 44464 0 1 20384
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1669390400
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_392
timestamp 1669390400
transform 1 0 45248 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_22_456
timestamp 1669390400
transform 1 0 52416 0 1 20384
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_460
timestamp 1669390400
transform 1 0 52864 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_463
timestamp 1669390400
transform 1 0 53200 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_22_527
timestamp 1669390400
transform 1 0 60368 0 1 20384
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_531
timestamp 1669390400
transform 1 0 60816 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_534
timestamp 1669390400
transform 1 0 61152 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_22_598
timestamp 1669390400
transform 1 0 68320 0 1 20384
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_602
timestamp 1669390400
transform 1 0 68768 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_605
timestamp 1669390400
transform 1 0 69104 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_22_669
timestamp 1669390400
transform 1 0 76272 0 1 20384
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_673
timestamp 1669390400
transform 1 0 76720 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_22_676
timestamp 1669390400
transform 1 0 77056 0 1 20384
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_22_684
timestamp 1669390400
transform 1 0 77952 0 1 20384
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_2
timestamp 1669390400
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_23_66
timestamp 1669390400
transform 1 0 8736 0 -1 21952
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1669390400
transform 1 0 9184 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1669390400
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_23_137
timestamp 1669390400
transform 1 0 16688 0 -1 21952
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1669390400
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_144
timestamp 1669390400
transform 1 0 17472 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_23_208
timestamp 1669390400
transform 1 0 24640 0 -1 21952
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1669390400
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1669390400
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_23_279
timestamp 1669390400
transform 1 0 32592 0 -1 21952
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1669390400
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1669390400
transform 1 0 33376 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_23_350
timestamp 1669390400
transform 1 0 40544 0 -1 21952
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1669390400
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_357
timestamp 1669390400
transform 1 0 41328 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_23_421
timestamp 1669390400
transform 1 0 48496 0 -1 21952
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_425
timestamp 1669390400
transform 1 0 48944 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_428
timestamp 1669390400
transform 1 0 49280 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_23_492
timestamp 1669390400
transform 1 0 56448 0 -1 21952
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_496
timestamp 1669390400
transform 1 0 56896 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_499
timestamp 1669390400
transform 1 0 57232 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_23_563
timestamp 1669390400
transform 1 0 64400 0 -1 21952
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_567
timestamp 1669390400
transform 1 0 64848 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_570
timestamp 1669390400
transform 1 0 65184 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_23_634
timestamp 1669390400
transform 1 0 72352 0 -1 21952
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_638
timestamp 1669390400
transform 1 0 72800 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_23_641
timestamp 1669390400
transform 1 0 73136 0 -1 21952
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_23_673
timestamp 1669390400
transform 1 0 76720 0 -1 21952
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_23_681
timestamp 1669390400
transform 1 0 77616 0 -1 21952
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_685
timestamp 1669390400
transform 1 0 78064 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_687
timestamp 1669390400
transform 1 0 78288 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_24_2
timestamp 1669390400
transform 1 0 1568 0 1 21952
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1669390400
transform 1 0 5152 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1669390400
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_24_101
timestamp 1669390400
transform 1 0 12656 0 1 21952
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1669390400
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1669390400
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_24_172
timestamp 1669390400
transform 1 0 20608 0 1 21952
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1669390400
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_179
timestamp 1669390400
transform 1 0 21392 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_24_243
timestamp 1669390400
transform 1 0 28560 0 1 21952
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1669390400
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1669390400
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_24_314
timestamp 1669390400
transform 1 0 36512 0 1 21952
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1669390400
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_321
timestamp 1669390400
transform 1 0 37296 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_24_385
timestamp 1669390400
transform 1 0 44464 0 1 21952
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1669390400
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_392
timestamp 1669390400
transform 1 0 45248 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_24_456
timestamp 1669390400
transform 1 0 52416 0 1 21952
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_460
timestamp 1669390400
transform 1 0 52864 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_463
timestamp 1669390400
transform 1 0 53200 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_24_527
timestamp 1669390400
transform 1 0 60368 0 1 21952
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_531
timestamp 1669390400
transform 1 0 60816 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_534
timestamp 1669390400
transform 1 0 61152 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_24_598
timestamp 1669390400
transform 1 0 68320 0 1 21952
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_602
timestamp 1669390400
transform 1 0 68768 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_605
timestamp 1669390400
transform 1 0 69104 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_24_669
timestamp 1669390400
transform 1 0 76272 0 1 21952
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_673
timestamp 1669390400
transform 1 0 76720 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_24_676
timestamp 1669390400
transform 1 0 77056 0 1 21952
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_24_684
timestamp 1669390400
transform 1 0 77952 0 1 21952
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_2
timestamp 1669390400
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_25_66
timestamp 1669390400
transform 1 0 8736 0 -1 23520
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1669390400
transform 1 0 9184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1669390400
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_25_137
timestamp 1669390400
transform 1 0 16688 0 -1 23520
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1669390400
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1669390400
transform 1 0 17472 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_25_208
timestamp 1669390400
transform 1 0 24640 0 -1 23520
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1669390400
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1669390400
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_25_279
timestamp 1669390400
transform 1 0 32592 0 -1 23520
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1669390400
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_286
timestamp 1669390400
transform 1 0 33376 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_25_350
timestamp 1669390400
transform 1 0 40544 0 -1 23520
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1669390400
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_357
timestamp 1669390400
transform 1 0 41328 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_25_421
timestamp 1669390400
transform 1 0 48496 0 -1 23520
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_425
timestamp 1669390400
transform 1 0 48944 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_428
timestamp 1669390400
transform 1 0 49280 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_25_492
timestamp 1669390400
transform 1 0 56448 0 -1 23520
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_496
timestamp 1669390400
transform 1 0 56896 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_499
timestamp 1669390400
transform 1 0 57232 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_25_563
timestamp 1669390400
transform 1 0 64400 0 -1 23520
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_567
timestamp 1669390400
transform 1 0 64848 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_570
timestamp 1669390400
transform 1 0 65184 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_25_634
timestamp 1669390400
transform 1 0 72352 0 -1 23520
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_638
timestamp 1669390400
transform 1 0 72800 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_25_641
timestamp 1669390400
transform 1 0 73136 0 -1 23520
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_25_673
timestamp 1669390400
transform 1 0 76720 0 -1 23520
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_25_681
timestamp 1669390400
transform 1 0 77616 0 -1 23520
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_685
timestamp 1669390400
transform 1 0 78064 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_687
timestamp 1669390400
transform 1 0 78288 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_26_2
timestamp 1669390400
transform 1 0 1568 0 1 23520
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1669390400
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1669390400
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_26_101
timestamp 1669390400
transform 1 0 12656 0 1 23520
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1669390400
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1669390400
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_26_172
timestamp 1669390400
transform 1 0 20608 0 1 23520
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1669390400
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_179
timestamp 1669390400
transform 1 0 21392 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_26_243
timestamp 1669390400
transform 1 0 28560 0 1 23520
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1669390400
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1669390400
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_26_314
timestamp 1669390400
transform 1 0 36512 0 1 23520
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1669390400
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_321
timestamp 1669390400
transform 1 0 37296 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_26_385
timestamp 1669390400
transform 1 0 44464 0 1 23520
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1669390400
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_392
timestamp 1669390400
transform 1 0 45248 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_26_456
timestamp 1669390400
transform 1 0 52416 0 1 23520
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_460
timestamp 1669390400
transform 1 0 52864 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_463
timestamp 1669390400
transform 1 0 53200 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_26_527
timestamp 1669390400
transform 1 0 60368 0 1 23520
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_531
timestamp 1669390400
transform 1 0 60816 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_534
timestamp 1669390400
transform 1 0 61152 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_26_598
timestamp 1669390400
transform 1 0 68320 0 1 23520
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_602
timestamp 1669390400
transform 1 0 68768 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_605
timestamp 1669390400
transform 1 0 69104 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_26_669
timestamp 1669390400
transform 1 0 76272 0 1 23520
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_673
timestamp 1669390400
transform 1 0 76720 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_26_676
timestamp 1669390400
transform 1 0 77056 0 1 23520
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_26_684
timestamp 1669390400
transform 1 0 77952 0 1 23520
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_2
timestamp 1669390400
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_27_66
timestamp 1669390400
transform 1 0 8736 0 -1 25088
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1669390400
transform 1 0 9184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1669390400
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_27_137
timestamp 1669390400
transform 1 0 16688 0 -1 25088
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1669390400
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1669390400
transform 1 0 17472 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_27_208
timestamp 1669390400
transform 1 0 24640 0 -1 25088
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1669390400
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_215
timestamp 1669390400
transform 1 0 25424 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_27_279
timestamp 1669390400
transform 1 0 32592 0 -1 25088
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1669390400
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1669390400
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_27_350
timestamp 1669390400
transform 1 0 40544 0 -1 25088
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1669390400
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_357
timestamp 1669390400
transform 1 0 41328 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_27_421
timestamp 1669390400
transform 1 0 48496 0 -1 25088
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_425
timestamp 1669390400
transform 1 0 48944 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_428
timestamp 1669390400
transform 1 0 49280 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_27_492
timestamp 1669390400
transform 1 0 56448 0 -1 25088
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_496
timestamp 1669390400
transform 1 0 56896 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_499
timestamp 1669390400
transform 1 0 57232 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_27_563
timestamp 1669390400
transform 1 0 64400 0 -1 25088
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_567
timestamp 1669390400
transform 1 0 64848 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_570
timestamp 1669390400
transform 1 0 65184 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_27_634
timestamp 1669390400
transform 1 0 72352 0 -1 25088
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_638
timestamp 1669390400
transform 1 0 72800 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_27_641
timestamp 1669390400
transform 1 0 73136 0 -1 25088
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_27_673
timestamp 1669390400
transform 1 0 76720 0 -1 25088
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_27_681
timestamp 1669390400
transform 1 0 77616 0 -1 25088
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_685
timestamp 1669390400
transform 1 0 78064 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_687
timestamp 1669390400
transform 1 0 78288 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_28_2
timestamp 1669390400
transform 1 0 1568 0 1 25088
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1669390400
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1669390400
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_28_101
timestamp 1669390400
transform 1 0 12656 0 1 25088
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1669390400
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1669390400
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_28_172
timestamp 1669390400
transform 1 0 20608 0 1 25088
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1669390400
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1669390400
transform 1 0 21392 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_28_243
timestamp 1669390400
transform 1 0 28560 0 1 25088
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1669390400
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1669390400
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_28_314
timestamp 1669390400
transform 1 0 36512 0 1 25088
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1669390400
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_321
timestamp 1669390400
transform 1 0 37296 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_28_385
timestamp 1669390400
transform 1 0 44464 0 1 25088
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1669390400
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_392
timestamp 1669390400
transform 1 0 45248 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_28_456
timestamp 1669390400
transform 1 0 52416 0 1 25088
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_460
timestamp 1669390400
transform 1 0 52864 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_463
timestamp 1669390400
transform 1 0 53200 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_28_527
timestamp 1669390400
transform 1 0 60368 0 1 25088
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_531
timestamp 1669390400
transform 1 0 60816 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_534
timestamp 1669390400
transform 1 0 61152 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_28_598
timestamp 1669390400
transform 1 0 68320 0 1 25088
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_602
timestamp 1669390400
transform 1 0 68768 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_605
timestamp 1669390400
transform 1 0 69104 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_28_669
timestamp 1669390400
transform 1 0 76272 0 1 25088
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_673
timestamp 1669390400
transform 1 0 76720 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_28_676
timestamp 1669390400
transform 1 0 77056 0 1 25088
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_28_684
timestamp 1669390400
transform 1 0 77952 0 1 25088
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1669390400
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_29_66
timestamp 1669390400
transform 1 0 8736 0 -1 26656
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1669390400
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1669390400
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_29_137
timestamp 1669390400
transform 1 0 16688 0 -1 26656
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1669390400
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1669390400
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_29_208
timestamp 1669390400
transform 1 0 24640 0 -1 26656
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1669390400
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1669390400
transform 1 0 25424 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_29_279
timestamp 1669390400
transform 1 0 32592 0 -1 26656
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1669390400
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1669390400
transform 1 0 33376 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_29_350
timestamp 1669390400
transform 1 0 40544 0 -1 26656
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1669390400
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_357
timestamp 1669390400
transform 1 0 41328 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_29_421
timestamp 1669390400
transform 1 0 48496 0 -1 26656
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_425
timestamp 1669390400
transform 1 0 48944 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_428
timestamp 1669390400
transform 1 0 49280 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_29_492
timestamp 1669390400
transform 1 0 56448 0 -1 26656
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_496
timestamp 1669390400
transform 1 0 56896 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_499
timestamp 1669390400
transform 1 0 57232 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_29_563
timestamp 1669390400
transform 1 0 64400 0 -1 26656
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_567
timestamp 1669390400
transform 1 0 64848 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_570
timestamp 1669390400
transform 1 0 65184 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_29_634
timestamp 1669390400
transform 1 0 72352 0 -1 26656
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_638
timestamp 1669390400
transform 1 0 72800 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_29_641
timestamp 1669390400
transform 1 0 73136 0 -1 26656
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_29_673
timestamp 1669390400
transform 1 0 76720 0 -1 26656
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_29_681
timestamp 1669390400
transform 1 0 77616 0 -1 26656
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_685
timestamp 1669390400
transform 1 0 78064 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_687
timestamp 1669390400
transform 1 0 78288 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_30_2
timestamp 1669390400
transform 1 0 1568 0 1 26656
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1669390400
transform 1 0 5152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1669390400
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_30_101
timestamp 1669390400
transform 1 0 12656 0 1 26656
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1669390400
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1669390400
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_30_172
timestamp 1669390400
transform 1 0 20608 0 1 26656
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1669390400
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1669390400
transform 1 0 21392 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_30_243
timestamp 1669390400
transform 1 0 28560 0 1 26656
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1669390400
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1669390400
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_30_314
timestamp 1669390400
transform 1 0 36512 0 1 26656
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1669390400
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_321
timestamp 1669390400
transform 1 0 37296 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_30_385
timestamp 1669390400
transform 1 0 44464 0 1 26656
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1669390400
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_392
timestamp 1669390400
transform 1 0 45248 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_30_456
timestamp 1669390400
transform 1 0 52416 0 1 26656
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_460
timestamp 1669390400
transform 1 0 52864 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_463
timestamp 1669390400
transform 1 0 53200 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_30_527
timestamp 1669390400
transform 1 0 60368 0 1 26656
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_531
timestamp 1669390400
transform 1 0 60816 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_534
timestamp 1669390400
transform 1 0 61152 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_30_598
timestamp 1669390400
transform 1 0 68320 0 1 26656
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_602
timestamp 1669390400
transform 1 0 68768 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_605
timestamp 1669390400
transform 1 0 69104 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_30_669
timestamp 1669390400
transform 1 0 76272 0 1 26656
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_673
timestamp 1669390400
transform 1 0 76720 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_30_676
timestamp 1669390400
transform 1 0 77056 0 1 26656
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_30_684
timestamp 1669390400
transform 1 0 77952 0 1 26656
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_2
timestamp 1669390400
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_31_66
timestamp 1669390400
transform 1 0 8736 0 -1 28224
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1669390400
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1669390400
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_31_137
timestamp 1669390400
transform 1 0 16688 0 -1 28224
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1669390400
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1669390400
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_31_208
timestamp 1669390400
transform 1 0 24640 0 -1 28224
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1669390400
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1669390400
transform 1 0 25424 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_31_279
timestamp 1669390400
transform 1 0 32592 0 -1 28224
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1669390400
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1669390400
transform 1 0 33376 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_31_350
timestamp 1669390400
transform 1 0 40544 0 -1 28224
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1669390400
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_357
timestamp 1669390400
transform 1 0 41328 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_31_421
timestamp 1669390400
transform 1 0 48496 0 -1 28224
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_425
timestamp 1669390400
transform 1 0 48944 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_428
timestamp 1669390400
transform 1 0 49280 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_31_492
timestamp 1669390400
transform 1 0 56448 0 -1 28224
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_496
timestamp 1669390400
transform 1 0 56896 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_499
timestamp 1669390400
transform 1 0 57232 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_31_563
timestamp 1669390400
transform 1 0 64400 0 -1 28224
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_567
timestamp 1669390400
transform 1 0 64848 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_570
timestamp 1669390400
transform 1 0 65184 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_31_634
timestamp 1669390400
transform 1 0 72352 0 -1 28224
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_638
timestamp 1669390400
transform 1 0 72800 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_31_641
timestamp 1669390400
transform 1 0 73136 0 -1 28224
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_31_673
timestamp 1669390400
transform 1 0 76720 0 -1 28224
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_31_681
timestamp 1669390400
transform 1 0 77616 0 -1 28224
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_685
timestamp 1669390400
transform 1 0 78064 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_687
timestamp 1669390400
transform 1 0 78288 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_32_2
timestamp 1669390400
transform 1 0 1568 0 1 28224
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1669390400
transform 1 0 5152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1669390400
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_32_101
timestamp 1669390400
transform 1 0 12656 0 1 28224
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1669390400
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1669390400
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_32_172
timestamp 1669390400
transform 1 0 20608 0 1 28224
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1669390400
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_179
timestamp 1669390400
transform 1 0 21392 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_32_243
timestamp 1669390400
transform 1 0 28560 0 1 28224
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1669390400
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1669390400
transform 1 0 29344 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_32_314
timestamp 1669390400
transform 1 0 36512 0 1 28224
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1669390400
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_321
timestamp 1669390400
transform 1 0 37296 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_32_385
timestamp 1669390400
transform 1 0 44464 0 1 28224
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1669390400
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_392
timestamp 1669390400
transform 1 0 45248 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_32_456
timestamp 1669390400
transform 1 0 52416 0 1 28224
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_460
timestamp 1669390400
transform 1 0 52864 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_463
timestamp 1669390400
transform 1 0 53200 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_32_527
timestamp 1669390400
transform 1 0 60368 0 1 28224
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_531
timestamp 1669390400
transform 1 0 60816 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_534
timestamp 1669390400
transform 1 0 61152 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_32_598
timestamp 1669390400
transform 1 0 68320 0 1 28224
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_602
timestamp 1669390400
transform 1 0 68768 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_605
timestamp 1669390400
transform 1 0 69104 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_32_669
timestamp 1669390400
transform 1 0 76272 0 1 28224
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_673
timestamp 1669390400
transform 1 0 76720 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_32_676
timestamp 1669390400
transform 1 0 77056 0 1 28224
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_32_684
timestamp 1669390400
transform 1 0 77952 0 1 28224
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1669390400
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_33_66
timestamp 1669390400
transform 1 0 8736 0 -1 29792
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1669390400
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1669390400
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_33_137
timestamp 1669390400
transform 1 0 16688 0 -1 29792
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1669390400
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1669390400
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_33_208
timestamp 1669390400
transform 1 0 24640 0 -1 29792
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1669390400
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1669390400
transform 1 0 25424 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_33_279
timestamp 1669390400
transform 1 0 32592 0 -1 29792
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1669390400
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1669390400
transform 1 0 33376 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_33_350
timestamp 1669390400
transform 1 0 40544 0 -1 29792
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1669390400
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_357
timestamp 1669390400
transform 1 0 41328 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_33_421
timestamp 1669390400
transform 1 0 48496 0 -1 29792
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_425
timestamp 1669390400
transform 1 0 48944 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_428
timestamp 1669390400
transform 1 0 49280 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_33_492
timestamp 1669390400
transform 1 0 56448 0 -1 29792
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_496
timestamp 1669390400
transform 1 0 56896 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_499
timestamp 1669390400
transform 1 0 57232 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_33_563
timestamp 1669390400
transform 1 0 64400 0 -1 29792
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_567
timestamp 1669390400
transform 1 0 64848 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_570
timestamp 1669390400
transform 1 0 65184 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_33_634
timestamp 1669390400
transform 1 0 72352 0 -1 29792
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_638
timestamp 1669390400
transform 1 0 72800 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_33_641
timestamp 1669390400
transform 1 0 73136 0 -1 29792
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_33_673
timestamp 1669390400
transform 1 0 76720 0 -1 29792
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_33_681
timestamp 1669390400
transform 1 0 77616 0 -1 29792
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_685
timestamp 1669390400
transform 1 0 78064 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_687
timestamp 1669390400
transform 1 0 78288 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_34_2
timestamp 1669390400
transform 1 0 1568 0 1 29792
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1669390400
transform 1 0 5152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1669390400
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_34_101
timestamp 1669390400
transform 1 0 12656 0 1 29792
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1669390400
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1669390400
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_34_172
timestamp 1669390400
transform 1 0 20608 0 1 29792
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1669390400
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1669390400
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_34_243
timestamp 1669390400
transform 1 0 28560 0 1 29792
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1669390400
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1669390400
transform 1 0 29344 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_34_314
timestamp 1669390400
transform 1 0 36512 0 1 29792
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1669390400
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_321
timestamp 1669390400
transform 1 0 37296 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_34_385
timestamp 1669390400
transform 1 0 44464 0 1 29792
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1669390400
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_392
timestamp 1669390400
transform 1 0 45248 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_34_456
timestamp 1669390400
transform 1 0 52416 0 1 29792
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_460
timestamp 1669390400
transform 1 0 52864 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_463
timestamp 1669390400
transform 1 0 53200 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_34_527
timestamp 1669390400
transform 1 0 60368 0 1 29792
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_531
timestamp 1669390400
transform 1 0 60816 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_534
timestamp 1669390400
transform 1 0 61152 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_34_598
timestamp 1669390400
transform 1 0 68320 0 1 29792
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_602
timestamp 1669390400
transform 1 0 68768 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_605
timestamp 1669390400
transform 1 0 69104 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_34_669
timestamp 1669390400
transform 1 0 76272 0 1 29792
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_673
timestamp 1669390400
transform 1 0 76720 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_34_676
timestamp 1669390400
transform 1 0 77056 0 1 29792
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_34_684
timestamp 1669390400
transform 1 0 77952 0 1 29792
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1669390400
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_35_66
timestamp 1669390400
transform 1 0 8736 0 -1 31360
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1669390400
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1669390400
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_35_137
timestamp 1669390400
transform 1 0 16688 0 -1 31360
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1669390400
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1669390400
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_35_208
timestamp 1669390400
transform 1 0 24640 0 -1 31360
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1669390400
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_215
timestamp 1669390400
transform 1 0 25424 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_35_279
timestamp 1669390400
transform 1 0 32592 0 -1 31360
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1669390400
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1669390400
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_35_350
timestamp 1669390400
transform 1 0 40544 0 -1 31360
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1669390400
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_357
timestamp 1669390400
transform 1 0 41328 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_35_421
timestamp 1669390400
transform 1 0 48496 0 -1 31360
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_425
timestamp 1669390400
transform 1 0 48944 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_428
timestamp 1669390400
transform 1 0 49280 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_35_492
timestamp 1669390400
transform 1 0 56448 0 -1 31360
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1669390400
transform 1 0 56896 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_499
timestamp 1669390400
transform 1 0 57232 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_35_563
timestamp 1669390400
transform 1 0 64400 0 -1 31360
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_567
timestamp 1669390400
transform 1 0 64848 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_570
timestamp 1669390400
transform 1 0 65184 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_35_634
timestamp 1669390400
transform 1 0 72352 0 -1 31360
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_638
timestamp 1669390400
transform 1 0 72800 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_35_641
timestamp 1669390400
transform 1 0 73136 0 -1 31360
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_35_673
timestamp 1669390400
transform 1 0 76720 0 -1 31360
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_35_681
timestamp 1669390400
transform 1 0 77616 0 -1 31360
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_685
timestamp 1669390400
transform 1 0 78064 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_687
timestamp 1669390400
transform 1 0 78288 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_36_2
timestamp 1669390400
transform 1 0 1568 0 1 31360
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1669390400
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1669390400
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_36_101
timestamp 1669390400
transform 1 0 12656 0 1 31360
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1669390400
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1669390400
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_36_172
timestamp 1669390400
transform 1 0 20608 0 1 31360
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1669390400
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1669390400
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_36_243
timestamp 1669390400
transform 1 0 28560 0 1 31360
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1669390400
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_250
timestamp 1669390400
transform 1 0 29344 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_36_314
timestamp 1669390400
transform 1 0 36512 0 1 31360
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1669390400
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_321
timestamp 1669390400
transform 1 0 37296 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_36_385
timestamp 1669390400
transform 1 0 44464 0 1 31360
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1669390400
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_392
timestamp 1669390400
transform 1 0 45248 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_36_456
timestamp 1669390400
transform 1 0 52416 0 1 31360
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1669390400
transform 1 0 52864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_463
timestamp 1669390400
transform 1 0 53200 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_36_527
timestamp 1669390400
transform 1 0 60368 0 1 31360
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_531
timestamp 1669390400
transform 1 0 60816 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_534
timestamp 1669390400
transform 1 0 61152 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_36_598
timestamp 1669390400
transform 1 0 68320 0 1 31360
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_602
timestamp 1669390400
transform 1 0 68768 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_605
timestamp 1669390400
transform 1 0 69104 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_36_669
timestamp 1669390400
transform 1 0 76272 0 1 31360
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_673
timestamp 1669390400
transform 1 0 76720 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_36_676
timestamp 1669390400
transform 1 0 77056 0 1 31360
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_36_684
timestamp 1669390400
transform 1 0 77952 0 1 31360
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1669390400
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_37_66
timestamp 1669390400
transform 1 0 8736 0 -1 32928
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1669390400
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1669390400
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_37_137
timestamp 1669390400
transform 1 0 16688 0 -1 32928
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1669390400
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1669390400
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_37_208
timestamp 1669390400
transform 1 0 24640 0 -1 32928
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1669390400
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_215
timestamp 1669390400
transform 1 0 25424 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_37_279
timestamp 1669390400
transform 1 0 32592 0 -1 32928
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1669390400
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_286
timestamp 1669390400
transform 1 0 33376 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_37_350
timestamp 1669390400
transform 1 0 40544 0 -1 32928
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1669390400
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_357
timestamp 1669390400
transform 1 0 41328 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_37_421
timestamp 1669390400
transform 1 0 48496 0 -1 32928
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_425
timestamp 1669390400
transform 1 0 48944 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_428
timestamp 1669390400
transform 1 0 49280 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_37_492
timestamp 1669390400
transform 1 0 56448 0 -1 32928
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_496
timestamp 1669390400
transform 1 0 56896 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_499
timestamp 1669390400
transform 1 0 57232 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_37_563
timestamp 1669390400
transform 1 0 64400 0 -1 32928
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_567
timestamp 1669390400
transform 1 0 64848 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_570
timestamp 1669390400
transform 1 0 65184 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_37_634
timestamp 1669390400
transform 1 0 72352 0 -1 32928
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_638
timestamp 1669390400
transform 1 0 72800 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_37_641
timestamp 1669390400
transform 1 0 73136 0 -1 32928
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_37_673
timestamp 1669390400
transform 1 0 76720 0 -1 32928
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_37_681
timestamp 1669390400
transform 1 0 77616 0 -1 32928
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_685
timestamp 1669390400
transform 1 0 78064 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_687
timestamp 1669390400
transform 1 0 78288 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_38_2
timestamp 1669390400
transform 1 0 1568 0 1 32928
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1669390400
transform 1 0 5152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1669390400
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_38_101
timestamp 1669390400
transform 1 0 12656 0 1 32928
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1669390400
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_108
timestamp 1669390400
transform 1 0 13440 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_38_172
timestamp 1669390400
transform 1 0 20608 0 1 32928
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1669390400
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1669390400
transform 1 0 21392 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_38_243
timestamp 1669390400
transform 1 0 28560 0 1 32928
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1669390400
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_250
timestamp 1669390400
transform 1 0 29344 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_38_314
timestamp 1669390400
transform 1 0 36512 0 1 32928
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1669390400
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_321
timestamp 1669390400
transform 1 0 37296 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_38_385
timestamp 1669390400
transform 1 0 44464 0 1 32928
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1669390400
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_392
timestamp 1669390400
transform 1 0 45248 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_38_456
timestamp 1669390400
transform 1 0 52416 0 1 32928
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_460
timestamp 1669390400
transform 1 0 52864 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_463
timestamp 1669390400
transform 1 0 53200 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_38_527
timestamp 1669390400
transform 1 0 60368 0 1 32928
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_531
timestamp 1669390400
transform 1 0 60816 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_534
timestamp 1669390400
transform 1 0 61152 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_38_598
timestamp 1669390400
transform 1 0 68320 0 1 32928
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_602
timestamp 1669390400
transform 1 0 68768 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_605
timestamp 1669390400
transform 1 0 69104 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_38_669
timestamp 1669390400
transform 1 0 76272 0 1 32928
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_673
timestamp 1669390400
transform 1 0 76720 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_38_676
timestamp 1669390400
transform 1 0 77056 0 1 32928
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_38_684
timestamp 1669390400
transform 1 0 77952 0 1 32928
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1669390400
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_39_66
timestamp 1669390400
transform 1 0 8736 0 -1 34496
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1669390400
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1669390400
transform 1 0 9520 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_39_137
timestamp 1669390400
transform 1 0 16688 0 -1 34496
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1669390400
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_144
timestamp 1669390400
transform 1 0 17472 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_39_208
timestamp 1669390400
transform 1 0 24640 0 -1 34496
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1669390400
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_215
timestamp 1669390400
transform 1 0 25424 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_39_279
timestamp 1669390400
transform 1 0 32592 0 -1 34496
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1669390400
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_286
timestamp 1669390400
transform 1 0 33376 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_39_350
timestamp 1669390400
transform 1 0 40544 0 -1 34496
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1669390400
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_357
timestamp 1669390400
transform 1 0 41328 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_39_421
timestamp 1669390400
transform 1 0 48496 0 -1 34496
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_425
timestamp 1669390400
transform 1 0 48944 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_428
timestamp 1669390400
transform 1 0 49280 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_39_492
timestamp 1669390400
transform 1 0 56448 0 -1 34496
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_496
timestamp 1669390400
transform 1 0 56896 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_499
timestamp 1669390400
transform 1 0 57232 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_39_563
timestamp 1669390400
transform 1 0 64400 0 -1 34496
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_567
timestamp 1669390400
transform 1 0 64848 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_570
timestamp 1669390400
transform 1 0 65184 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_39_634
timestamp 1669390400
transform 1 0 72352 0 -1 34496
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_638
timestamp 1669390400
transform 1 0 72800 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_39_641
timestamp 1669390400
transform 1 0 73136 0 -1 34496
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_39_673
timestamp 1669390400
transform 1 0 76720 0 -1 34496
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_39_681
timestamp 1669390400
transform 1 0 77616 0 -1 34496
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_685
timestamp 1669390400
transform 1 0 78064 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_687
timestamp 1669390400
transform 1 0 78288 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_40_2
timestamp 1669390400
transform 1 0 1568 0 1 34496
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1669390400
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1669390400
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_40_101
timestamp 1669390400
transform 1 0 12656 0 1 34496
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1669390400
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_108
timestamp 1669390400
transform 1 0 13440 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_40_172
timestamp 1669390400
transform 1 0 20608 0 1 34496
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1669390400
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_179
timestamp 1669390400
transform 1 0 21392 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_40_243
timestamp 1669390400
transform 1 0 28560 0 1 34496
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1669390400
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_250
timestamp 1669390400
transform 1 0 29344 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_40_314
timestamp 1669390400
transform 1 0 36512 0 1 34496
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1669390400
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_321
timestamp 1669390400
transform 1 0 37296 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_40_385
timestamp 1669390400
transform 1 0 44464 0 1 34496
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1669390400
transform 1 0 44912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_392
timestamp 1669390400
transform 1 0 45248 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_40_456
timestamp 1669390400
transform 1 0 52416 0 1 34496
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_460
timestamp 1669390400
transform 1 0 52864 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_463
timestamp 1669390400
transform 1 0 53200 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_40_527
timestamp 1669390400
transform 1 0 60368 0 1 34496
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_531
timestamp 1669390400
transform 1 0 60816 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_534
timestamp 1669390400
transform 1 0 61152 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_40_598
timestamp 1669390400
transform 1 0 68320 0 1 34496
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_602
timestamp 1669390400
transform 1 0 68768 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_605
timestamp 1669390400
transform 1 0 69104 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_40_669
timestamp 1669390400
transform 1 0 76272 0 1 34496
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_673
timestamp 1669390400
transform 1 0 76720 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_40_676
timestamp 1669390400
transform 1 0 77056 0 1 34496
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_40_684
timestamp 1669390400
transform 1 0 77952 0 1 34496
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_2
timestamp 1669390400
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_41_66
timestamp 1669390400
transform 1 0 8736 0 -1 36064
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1669390400
transform 1 0 9184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1669390400
transform 1 0 9520 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_41_137
timestamp 1669390400
transform 1 0 16688 0 -1 36064
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1669390400
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_144
timestamp 1669390400
transform 1 0 17472 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_41_208
timestamp 1669390400
transform 1 0 24640 0 -1 36064
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1669390400
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1669390400
transform 1 0 25424 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_41_279
timestamp 1669390400
transform 1 0 32592 0 -1 36064
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1669390400
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_286
timestamp 1669390400
transform 1 0 33376 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_41_350
timestamp 1669390400
transform 1 0 40544 0 -1 36064
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1669390400
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_357
timestamp 1669390400
transform 1 0 41328 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_41_421
timestamp 1669390400
transform 1 0 48496 0 -1 36064
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_425
timestamp 1669390400
transform 1 0 48944 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_428
timestamp 1669390400
transform 1 0 49280 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_41_492
timestamp 1669390400
transform 1 0 56448 0 -1 36064
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_496
timestamp 1669390400
transform 1 0 56896 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_499
timestamp 1669390400
transform 1 0 57232 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_41_563
timestamp 1669390400
transform 1 0 64400 0 -1 36064
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_567
timestamp 1669390400
transform 1 0 64848 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_570
timestamp 1669390400
transform 1 0 65184 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_41_634
timestamp 1669390400
transform 1 0 72352 0 -1 36064
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_638
timestamp 1669390400
transform 1 0 72800 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_41_641
timestamp 1669390400
transform 1 0 73136 0 -1 36064
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_41_673
timestamp 1669390400
transform 1 0 76720 0 -1 36064
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_41_681
timestamp 1669390400
transform 1 0 77616 0 -1 36064
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_685
timestamp 1669390400
transform 1 0 78064 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_687
timestamp 1669390400
transform 1 0 78288 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_42_2
timestamp 1669390400
transform 1 0 1568 0 1 36064
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1669390400
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_37
timestamp 1669390400
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_42_101
timestamp 1669390400
transform 1 0 12656 0 1 36064
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1669390400
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_108
timestamp 1669390400
transform 1 0 13440 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_42_172
timestamp 1669390400
transform 1 0 20608 0 1 36064
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_176
timestamp 1669390400
transform 1 0 21056 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_179
timestamp 1669390400
transform 1 0 21392 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_42_243
timestamp 1669390400
transform 1 0 28560 0 1 36064
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1669390400
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_250
timestamp 1669390400
transform 1 0 29344 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_42_314
timestamp 1669390400
transform 1 0 36512 0 1 36064
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_318
timestamp 1669390400
transform 1 0 36960 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_321
timestamp 1669390400
transform 1 0 37296 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_42_385
timestamp 1669390400
transform 1 0 44464 0 1 36064
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_389
timestamp 1669390400
transform 1 0 44912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_392
timestamp 1669390400
transform 1 0 45248 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_42_456
timestamp 1669390400
transform 1 0 52416 0 1 36064
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_460
timestamp 1669390400
transform 1 0 52864 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_463
timestamp 1669390400
transform 1 0 53200 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_42_527
timestamp 1669390400
transform 1 0 60368 0 1 36064
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_531
timestamp 1669390400
transform 1 0 60816 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_534
timestamp 1669390400
transform 1 0 61152 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_42_598
timestamp 1669390400
transform 1 0 68320 0 1 36064
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_602
timestamp 1669390400
transform 1 0 68768 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_605
timestamp 1669390400
transform 1 0 69104 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_42_669
timestamp 1669390400
transform 1 0 76272 0 1 36064
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_673
timestamp 1669390400
transform 1 0 76720 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_42_676
timestamp 1669390400
transform 1 0 77056 0 1 36064
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_42_684
timestamp 1669390400
transform 1 0 77952 0 1 36064
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_2
timestamp 1669390400
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_43_66
timestamp 1669390400
transform 1 0 8736 0 -1 37632
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_70
timestamp 1669390400
transform 1 0 9184 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_73
timestamp 1669390400
transform 1 0 9520 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_43_137
timestamp 1669390400
transform 1 0 16688 0 -1 37632
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1669390400
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_144
timestamp 1669390400
transform 1 0 17472 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_43_208
timestamp 1669390400
transform 1 0 24640 0 -1 37632
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1669390400
transform 1 0 25088 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_215
timestamp 1669390400
transform 1 0 25424 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_43_279
timestamp 1669390400
transform 1 0 32592 0 -1 37632
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1669390400
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_286
timestamp 1669390400
transform 1 0 33376 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_43_350
timestamp 1669390400
transform 1 0 40544 0 -1 37632
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_354
timestamp 1669390400
transform 1 0 40992 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_357
timestamp 1669390400
transform 1 0 41328 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_43_421
timestamp 1669390400
transform 1 0 48496 0 -1 37632
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_425
timestamp 1669390400
transform 1 0 48944 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_428
timestamp 1669390400
transform 1 0 49280 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_43_492
timestamp 1669390400
transform 1 0 56448 0 -1 37632
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_496
timestamp 1669390400
transform 1 0 56896 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_499
timestamp 1669390400
transform 1 0 57232 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_43_563
timestamp 1669390400
transform 1 0 64400 0 -1 37632
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_567
timestamp 1669390400
transform 1 0 64848 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_570
timestamp 1669390400
transform 1 0 65184 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_43_634
timestamp 1669390400
transform 1 0 72352 0 -1 37632
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_638
timestamp 1669390400
transform 1 0 72800 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_43_641
timestamp 1669390400
transform 1 0 73136 0 -1 37632
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_43_673
timestamp 1669390400
transform 1 0 76720 0 -1 37632
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_43_681
timestamp 1669390400
transform 1 0 77616 0 -1 37632
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_685
timestamp 1669390400
transform 1 0 78064 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_687
timestamp 1669390400
transform 1 0 78288 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_44_2
timestamp 1669390400
transform 1 0 1568 0 1 37632
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_34
timestamp 1669390400
transform 1 0 5152 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_37
timestamp 1669390400
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_44_101
timestamp 1669390400
transform 1 0 12656 0 1 37632
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1669390400
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_108
timestamp 1669390400
transform 1 0 13440 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_44_172
timestamp 1669390400
transform 1 0 20608 0 1 37632
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1669390400
transform 1 0 21056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_179
timestamp 1669390400
transform 1 0 21392 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_44_243
timestamp 1669390400
transform 1 0 28560 0 1 37632
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_247
timestamp 1669390400
transform 1 0 29008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_250
timestamp 1669390400
transform 1 0 29344 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_44_314
timestamp 1669390400
transform 1 0 36512 0 1 37632
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_318
timestamp 1669390400
transform 1 0 36960 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_321
timestamp 1669390400
transform 1 0 37296 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_44_385
timestamp 1669390400
transform 1 0 44464 0 1 37632
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_389
timestamp 1669390400
transform 1 0 44912 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_392
timestamp 1669390400
transform 1 0 45248 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_44_456
timestamp 1669390400
transform 1 0 52416 0 1 37632
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_460
timestamp 1669390400
transform 1 0 52864 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_463
timestamp 1669390400
transform 1 0 53200 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_44_527
timestamp 1669390400
transform 1 0 60368 0 1 37632
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_531
timestamp 1669390400
transform 1 0 60816 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_534
timestamp 1669390400
transform 1 0 61152 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_44_598
timestamp 1669390400
transform 1 0 68320 0 1 37632
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_602
timestamp 1669390400
transform 1 0 68768 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_605
timestamp 1669390400
transform 1 0 69104 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_44_669
timestamp 1669390400
transform 1 0 76272 0 1 37632
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_673
timestamp 1669390400
transform 1 0 76720 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_44_676
timestamp 1669390400
transform 1 0 77056 0 1 37632
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_44_684
timestamp 1669390400
transform 1 0 77952 0 1 37632
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_2
timestamp 1669390400
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_45_66
timestamp 1669390400
transform 1 0 8736 0 -1 39200
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_70
timestamp 1669390400
transform 1 0 9184 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_73
timestamp 1669390400
transform 1 0 9520 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_45_137
timestamp 1669390400
transform 1 0 16688 0 -1 39200
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1669390400
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_144
timestamp 1669390400
transform 1 0 17472 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_45_208
timestamp 1669390400
transform 1 0 24640 0 -1 39200
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1669390400
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_215
timestamp 1669390400
transform 1 0 25424 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_45_279
timestamp 1669390400
transform 1 0 32592 0 -1 39200
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1669390400
transform 1 0 33040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_286
timestamp 1669390400
transform 1 0 33376 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_45_350
timestamp 1669390400
transform 1 0 40544 0 -1 39200
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_354
timestamp 1669390400
transform 1 0 40992 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_357
timestamp 1669390400
transform 1 0 41328 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_45_421
timestamp 1669390400
transform 1 0 48496 0 -1 39200
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_425
timestamp 1669390400
transform 1 0 48944 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_428
timestamp 1669390400
transform 1 0 49280 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_45_492
timestamp 1669390400
transform 1 0 56448 0 -1 39200
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_496
timestamp 1669390400
transform 1 0 56896 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_499
timestamp 1669390400
transform 1 0 57232 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_45_563
timestamp 1669390400
transform 1 0 64400 0 -1 39200
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_567
timestamp 1669390400
transform 1 0 64848 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_570
timestamp 1669390400
transform 1 0 65184 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_45_634
timestamp 1669390400
transform 1 0 72352 0 -1 39200
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_638
timestamp 1669390400
transform 1 0 72800 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_45_641
timestamp 1669390400
transform 1 0 73136 0 -1 39200
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_45_673
timestamp 1669390400
transform 1 0 76720 0 -1 39200
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_45_681
timestamp 1669390400
transform 1 0 77616 0 -1 39200
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_685
timestamp 1669390400
transform 1 0 78064 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_687
timestamp 1669390400
transform 1 0 78288 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_46_2
timestamp 1669390400
transform 1 0 1568 0 1 39200
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1669390400
transform 1 0 5152 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_37
timestamp 1669390400
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_46_101
timestamp 1669390400
transform 1 0 12656 0 1 39200
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1669390400
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_108
timestamp 1669390400
transform 1 0 13440 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_46_172
timestamp 1669390400
transform 1 0 20608 0 1 39200
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1669390400
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_179
timestamp 1669390400
transform 1 0 21392 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_46_243
timestamp 1669390400
transform 1 0 28560 0 1 39200
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1669390400
transform 1 0 29008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_250
timestamp 1669390400
transform 1 0 29344 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_46_314
timestamp 1669390400
transform 1 0 36512 0 1 39200
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_318
timestamp 1669390400
transform 1 0 36960 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_321
timestamp 1669390400
transform 1 0 37296 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_46_385
timestamp 1669390400
transform 1 0 44464 0 1 39200
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_389
timestamp 1669390400
transform 1 0 44912 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_392
timestamp 1669390400
transform 1 0 45248 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_46_456
timestamp 1669390400
transform 1 0 52416 0 1 39200
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_460
timestamp 1669390400
transform 1 0 52864 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_463
timestamp 1669390400
transform 1 0 53200 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_46_527
timestamp 1669390400
transform 1 0 60368 0 1 39200
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_531
timestamp 1669390400
transform 1 0 60816 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_534
timestamp 1669390400
transform 1 0 61152 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_46_598
timestamp 1669390400
transform 1 0 68320 0 1 39200
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_602
timestamp 1669390400
transform 1 0 68768 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_605
timestamp 1669390400
transform 1 0 69104 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_46_669
timestamp 1669390400
transform 1 0 76272 0 1 39200
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_673
timestamp 1669390400
transform 1 0 76720 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_46_676
timestamp 1669390400
transform 1 0 77056 0 1 39200
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_46_684
timestamp 1669390400
transform 1 0 77952 0 1 39200
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_2
timestamp 1669390400
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_47_66
timestamp 1669390400
transform 1 0 8736 0 -1 40768
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_70
timestamp 1669390400
transform 1 0 9184 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_73
timestamp 1669390400
transform 1 0 9520 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_47_137
timestamp 1669390400
transform 1 0 16688 0 -1 40768
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1669390400
transform 1 0 17136 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_144
timestamp 1669390400
transform 1 0 17472 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_47_208
timestamp 1669390400
transform 1 0 24640 0 -1 40768
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1669390400
transform 1 0 25088 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_215
timestamp 1669390400
transform 1 0 25424 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_47_279
timestamp 1669390400
transform 1 0 32592 0 -1 40768
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_283
timestamp 1669390400
transform 1 0 33040 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_286
timestamp 1669390400
transform 1 0 33376 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_47_350
timestamp 1669390400
transform 1 0 40544 0 -1 40768
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_354
timestamp 1669390400
transform 1 0 40992 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_357
timestamp 1669390400
transform 1 0 41328 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_47_421
timestamp 1669390400
transform 1 0 48496 0 -1 40768
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_425
timestamp 1669390400
transform 1 0 48944 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_428
timestamp 1669390400
transform 1 0 49280 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_47_492
timestamp 1669390400
transform 1 0 56448 0 -1 40768
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_496
timestamp 1669390400
transform 1 0 56896 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_499
timestamp 1669390400
transform 1 0 57232 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_47_563
timestamp 1669390400
transform 1 0 64400 0 -1 40768
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_567
timestamp 1669390400
transform 1 0 64848 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_570
timestamp 1669390400
transform 1 0 65184 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_47_634
timestamp 1669390400
transform 1 0 72352 0 -1 40768
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_638
timestamp 1669390400
transform 1 0 72800 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_47_641
timestamp 1669390400
transform 1 0 73136 0 -1 40768
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_47_673
timestamp 1669390400
transform 1 0 76720 0 -1 40768
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_47_681
timestamp 1669390400
transform 1 0 77616 0 -1 40768
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_685
timestamp 1669390400
transform 1 0 78064 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_687
timestamp 1669390400
transform 1 0 78288 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_48_2
timestamp 1669390400
transform 1 0 1568 0 1 40768
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_34
timestamp 1669390400
transform 1 0 5152 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_37
timestamp 1669390400
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_48_101
timestamp 1669390400
transform 1 0 12656 0 1 40768
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1669390400
transform 1 0 13104 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_108
timestamp 1669390400
transform 1 0 13440 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_48_172
timestamp 1669390400
transform 1 0 20608 0 1 40768
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1669390400
transform 1 0 21056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_179
timestamp 1669390400
transform 1 0 21392 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_48_243
timestamp 1669390400
transform 1 0 28560 0 1 40768
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_247
timestamp 1669390400
transform 1 0 29008 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_250
timestamp 1669390400
transform 1 0 29344 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_48_314
timestamp 1669390400
transform 1 0 36512 0 1 40768
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_318
timestamp 1669390400
transform 1 0 36960 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_321
timestamp 1669390400
transform 1 0 37296 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_48_385
timestamp 1669390400
transform 1 0 44464 0 1 40768
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_389
timestamp 1669390400
transform 1 0 44912 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_392
timestamp 1669390400
transform 1 0 45248 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_48_456
timestamp 1669390400
transform 1 0 52416 0 1 40768
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_460
timestamp 1669390400
transform 1 0 52864 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_463
timestamp 1669390400
transform 1 0 53200 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_48_527
timestamp 1669390400
transform 1 0 60368 0 1 40768
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_531
timestamp 1669390400
transform 1 0 60816 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_534
timestamp 1669390400
transform 1 0 61152 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_48_598
timestamp 1669390400
transform 1 0 68320 0 1 40768
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_602
timestamp 1669390400
transform 1 0 68768 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_605
timestamp 1669390400
transform 1 0 69104 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_48_669
timestamp 1669390400
transform 1 0 76272 0 1 40768
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_673
timestamp 1669390400
transform 1 0 76720 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_48_676
timestamp 1669390400
transform 1 0 77056 0 1 40768
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_48_684
timestamp 1669390400
transform 1 0 77952 0 1 40768
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_2
timestamp 1669390400
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_49_66
timestamp 1669390400
transform 1 0 8736 0 -1 42336
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_70
timestamp 1669390400
transform 1 0 9184 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_73
timestamp 1669390400
transform 1 0 9520 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_49_137
timestamp 1669390400
transform 1 0 16688 0 -1 42336
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1669390400
transform 1 0 17136 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_144
timestamp 1669390400
transform 1 0 17472 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_49_208
timestamp 1669390400
transform 1 0 24640 0 -1 42336
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1669390400
transform 1 0 25088 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_215
timestamp 1669390400
transform 1 0 25424 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_49_279
timestamp 1669390400
transform 1 0 32592 0 -1 42336
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_283
timestamp 1669390400
transform 1 0 33040 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_286
timestamp 1669390400
transform 1 0 33376 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_49_350
timestamp 1669390400
transform 1 0 40544 0 -1 42336
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_354
timestamp 1669390400
transform 1 0 40992 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_357
timestamp 1669390400
transform 1 0 41328 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_49_421
timestamp 1669390400
transform 1 0 48496 0 -1 42336
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_425
timestamp 1669390400
transform 1 0 48944 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_428
timestamp 1669390400
transform 1 0 49280 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_49_492
timestamp 1669390400
transform 1 0 56448 0 -1 42336
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_496
timestamp 1669390400
transform 1 0 56896 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_499
timestamp 1669390400
transform 1 0 57232 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_49_563
timestamp 1669390400
transform 1 0 64400 0 -1 42336
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_567
timestamp 1669390400
transform 1 0 64848 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_570
timestamp 1669390400
transform 1 0 65184 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_49_634
timestamp 1669390400
transform 1 0 72352 0 -1 42336
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_638
timestamp 1669390400
transform 1 0 72800 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_49_641
timestamp 1669390400
transform 1 0 73136 0 -1 42336
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_49_673
timestamp 1669390400
transform 1 0 76720 0 -1 42336
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_49_681
timestamp 1669390400
transform 1 0 77616 0 -1 42336
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_685
timestamp 1669390400
transform 1 0 78064 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_687
timestamp 1669390400
transform 1 0 78288 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_50_2
timestamp 1669390400
transform 1 0 1568 0 1 42336
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1669390400
transform 1 0 5152 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_37
timestamp 1669390400
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_50_101
timestamp 1669390400
transform 1 0 12656 0 1 42336
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1669390400
transform 1 0 13104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_108
timestamp 1669390400
transform 1 0 13440 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_50_172
timestamp 1669390400
transform 1 0 20608 0 1 42336
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_176
timestamp 1669390400
transform 1 0 21056 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_179
timestamp 1669390400
transform 1 0 21392 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_50_243
timestamp 1669390400
transform 1 0 28560 0 1 42336
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_247
timestamp 1669390400
transform 1 0 29008 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_250
timestamp 1669390400
transform 1 0 29344 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_50_314
timestamp 1669390400
transform 1 0 36512 0 1 42336
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_318
timestamp 1669390400
transform 1 0 36960 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_321
timestamp 1669390400
transform 1 0 37296 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_50_385
timestamp 1669390400
transform 1 0 44464 0 1 42336
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_389
timestamp 1669390400
transform 1 0 44912 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_392
timestamp 1669390400
transform 1 0 45248 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_50_456
timestamp 1669390400
transform 1 0 52416 0 1 42336
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_460
timestamp 1669390400
transform 1 0 52864 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_463
timestamp 1669390400
transform 1 0 53200 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_50_527
timestamp 1669390400
transform 1 0 60368 0 1 42336
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_531
timestamp 1669390400
transform 1 0 60816 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_534
timestamp 1669390400
transform 1 0 61152 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_50_598
timestamp 1669390400
transform 1 0 68320 0 1 42336
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_602
timestamp 1669390400
transform 1 0 68768 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_605
timestamp 1669390400
transform 1 0 69104 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_50_669
timestamp 1669390400
transform 1 0 76272 0 1 42336
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_673
timestamp 1669390400
transform 1 0 76720 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_50_676
timestamp 1669390400
transform 1 0 77056 0 1 42336
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_50_684
timestamp 1669390400
transform 1 0 77952 0 1 42336
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_2
timestamp 1669390400
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_51_66
timestamp 1669390400
transform 1 0 8736 0 -1 43904
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_70
timestamp 1669390400
transform 1 0 9184 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_73
timestamp 1669390400
transform 1 0 9520 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_51_137
timestamp 1669390400
transform 1 0 16688 0 -1 43904
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_141
timestamp 1669390400
transform 1 0 17136 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_144
timestamp 1669390400
transform 1 0 17472 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_51_208
timestamp 1669390400
transform 1 0 24640 0 -1 43904
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1669390400
transform 1 0 25088 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_215
timestamp 1669390400
transform 1 0 25424 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_51_279
timestamp 1669390400
transform 1 0 32592 0 -1 43904
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_283
timestamp 1669390400
transform 1 0 33040 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_286
timestamp 1669390400
transform 1 0 33376 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_51_350
timestamp 1669390400
transform 1 0 40544 0 -1 43904
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_354
timestamp 1669390400
transform 1 0 40992 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_357
timestamp 1669390400
transform 1 0 41328 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_51_421
timestamp 1669390400
transform 1 0 48496 0 -1 43904
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_425
timestamp 1669390400
transform 1 0 48944 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_428
timestamp 1669390400
transform 1 0 49280 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_51_492
timestamp 1669390400
transform 1 0 56448 0 -1 43904
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_496
timestamp 1669390400
transform 1 0 56896 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_499
timestamp 1669390400
transform 1 0 57232 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_51_563
timestamp 1669390400
transform 1 0 64400 0 -1 43904
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_567
timestamp 1669390400
transform 1 0 64848 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_570
timestamp 1669390400
transform 1 0 65184 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_51_634
timestamp 1669390400
transform 1 0 72352 0 -1 43904
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_638
timestamp 1669390400
transform 1 0 72800 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_51_641
timestamp 1669390400
transform 1 0 73136 0 -1 43904
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_51_673
timestamp 1669390400
transform 1 0 76720 0 -1 43904
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_51_681
timestamp 1669390400
transform 1 0 77616 0 -1 43904
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_685
timestamp 1669390400
transform 1 0 78064 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_687
timestamp 1669390400
transform 1 0 78288 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_52_2
timestamp 1669390400
transform 1 0 1568 0 1 43904
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_34
timestamp 1669390400
transform 1 0 5152 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_37
timestamp 1669390400
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_52_101
timestamp 1669390400
transform 1 0 12656 0 1 43904
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_105
timestamp 1669390400
transform 1 0 13104 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_108
timestamp 1669390400
transform 1 0 13440 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_52_172
timestamp 1669390400
transform 1 0 20608 0 1 43904
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1669390400
transform 1 0 21056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_179
timestamp 1669390400
transform 1 0 21392 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_52_243
timestamp 1669390400
transform 1 0 28560 0 1 43904
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_247
timestamp 1669390400
transform 1 0 29008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_250
timestamp 1669390400
transform 1 0 29344 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_52_314
timestamp 1669390400
transform 1 0 36512 0 1 43904
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_318
timestamp 1669390400
transform 1 0 36960 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_321
timestamp 1669390400
transform 1 0 37296 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_52_385
timestamp 1669390400
transform 1 0 44464 0 1 43904
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_389
timestamp 1669390400
transform 1 0 44912 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_392
timestamp 1669390400
transform 1 0 45248 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_52_456
timestamp 1669390400
transform 1 0 52416 0 1 43904
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_460
timestamp 1669390400
transform 1 0 52864 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_463
timestamp 1669390400
transform 1 0 53200 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_52_527
timestamp 1669390400
transform 1 0 60368 0 1 43904
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_531
timestamp 1669390400
transform 1 0 60816 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_534
timestamp 1669390400
transform 1 0 61152 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_52_598
timestamp 1669390400
transform 1 0 68320 0 1 43904
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_602
timestamp 1669390400
transform 1 0 68768 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_605
timestamp 1669390400
transform 1 0 69104 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_52_669
timestamp 1669390400
transform 1 0 76272 0 1 43904
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_673
timestamp 1669390400
transform 1 0 76720 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_52_676
timestamp 1669390400
transform 1 0 77056 0 1 43904
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_52_684
timestamp 1669390400
transform 1 0 77952 0 1 43904
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_2
timestamp 1669390400
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_53_66
timestamp 1669390400
transform 1 0 8736 0 -1 45472
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_70
timestamp 1669390400
transform 1 0 9184 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_73
timestamp 1669390400
transform 1 0 9520 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_53_137
timestamp 1669390400
transform 1 0 16688 0 -1 45472
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_141
timestamp 1669390400
transform 1 0 17136 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_144
timestamp 1669390400
transform 1 0 17472 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_53_208
timestamp 1669390400
transform 1 0 24640 0 -1 45472
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1669390400
transform 1 0 25088 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_215
timestamp 1669390400
transform 1 0 25424 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_53_279
timestamp 1669390400
transform 1 0 32592 0 -1 45472
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1669390400
transform 1 0 33040 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_286
timestamp 1669390400
transform 1 0 33376 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_53_350
timestamp 1669390400
transform 1 0 40544 0 -1 45472
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_354
timestamp 1669390400
transform 1 0 40992 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_357
timestamp 1669390400
transform 1 0 41328 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_53_421
timestamp 1669390400
transform 1 0 48496 0 -1 45472
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_425
timestamp 1669390400
transform 1 0 48944 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_428
timestamp 1669390400
transform 1 0 49280 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_53_492
timestamp 1669390400
transform 1 0 56448 0 -1 45472
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_496
timestamp 1669390400
transform 1 0 56896 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_499
timestamp 1669390400
transform 1 0 57232 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_53_563
timestamp 1669390400
transform 1 0 64400 0 -1 45472
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_567
timestamp 1669390400
transform 1 0 64848 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_570
timestamp 1669390400
transform 1 0 65184 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_53_634
timestamp 1669390400
transform 1 0 72352 0 -1 45472
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_638
timestamp 1669390400
transform 1 0 72800 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_53_641
timestamp 1669390400
transform 1 0 73136 0 -1 45472
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_53_673
timestamp 1669390400
transform 1 0 76720 0 -1 45472
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_53_681
timestamp 1669390400
transform 1 0 77616 0 -1 45472
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_685
timestamp 1669390400
transform 1 0 78064 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_687
timestamp 1669390400
transform 1 0 78288 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_54_2
timestamp 1669390400
transform 1 0 1568 0 1 45472
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_34
timestamp 1669390400
transform 1 0 5152 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_37
timestamp 1669390400
transform 1 0 5488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_54_101
timestamp 1669390400
transform 1 0 12656 0 1 45472
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_105
timestamp 1669390400
transform 1 0 13104 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_108
timestamp 1669390400
transform 1 0 13440 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_54_172
timestamp 1669390400
transform 1 0 20608 0 1 45472
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_176
timestamp 1669390400
transform 1 0 21056 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_179
timestamp 1669390400
transform 1 0 21392 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_54_243
timestamp 1669390400
transform 1 0 28560 0 1 45472
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_247
timestamp 1669390400
transform 1 0 29008 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_250
timestamp 1669390400
transform 1 0 29344 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_54_314
timestamp 1669390400
transform 1 0 36512 0 1 45472
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_318
timestamp 1669390400
transform 1 0 36960 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_321
timestamp 1669390400
transform 1 0 37296 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_54_385
timestamp 1669390400
transform 1 0 44464 0 1 45472
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_389
timestamp 1669390400
transform 1 0 44912 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_392
timestamp 1669390400
transform 1 0 45248 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_54_456
timestamp 1669390400
transform 1 0 52416 0 1 45472
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_460
timestamp 1669390400
transform 1 0 52864 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_463
timestamp 1669390400
transform 1 0 53200 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_54_527
timestamp 1669390400
transform 1 0 60368 0 1 45472
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_531
timestamp 1669390400
transform 1 0 60816 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_534
timestamp 1669390400
transform 1 0 61152 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_54_598
timestamp 1669390400
transform 1 0 68320 0 1 45472
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_602
timestamp 1669390400
transform 1 0 68768 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_605
timestamp 1669390400
transform 1 0 69104 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_54_669
timestamp 1669390400
transform 1 0 76272 0 1 45472
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_673
timestamp 1669390400
transform 1 0 76720 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_54_676
timestamp 1669390400
transform 1 0 77056 0 1 45472
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_54_684
timestamp 1669390400
transform 1 0 77952 0 1 45472
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_2
timestamp 1669390400
transform 1 0 1568 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_55_66
timestamp 1669390400
transform 1 0 8736 0 -1 47040
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_70
timestamp 1669390400
transform 1 0 9184 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_73
timestamp 1669390400
transform 1 0 9520 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_55_137
timestamp 1669390400
transform 1 0 16688 0 -1 47040
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_141
timestamp 1669390400
transform 1 0 17136 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_144
timestamp 1669390400
transform 1 0 17472 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_55_208
timestamp 1669390400
transform 1 0 24640 0 -1 47040
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_212
timestamp 1669390400
transform 1 0 25088 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_215
timestamp 1669390400
transform 1 0 25424 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_55_279
timestamp 1669390400
transform 1 0 32592 0 -1 47040
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_283
timestamp 1669390400
transform 1 0 33040 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_286
timestamp 1669390400
transform 1 0 33376 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_55_350
timestamp 1669390400
transform 1 0 40544 0 -1 47040
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_354
timestamp 1669390400
transform 1 0 40992 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_357
timestamp 1669390400
transform 1 0 41328 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_55_421
timestamp 1669390400
transform 1 0 48496 0 -1 47040
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_425
timestamp 1669390400
transform 1 0 48944 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_428
timestamp 1669390400
transform 1 0 49280 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_55_492
timestamp 1669390400
transform 1 0 56448 0 -1 47040
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_496
timestamp 1669390400
transform 1 0 56896 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_499
timestamp 1669390400
transform 1 0 57232 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_55_563
timestamp 1669390400
transform 1 0 64400 0 -1 47040
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_567
timestamp 1669390400
transform 1 0 64848 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_570
timestamp 1669390400
transform 1 0 65184 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_55_634
timestamp 1669390400
transform 1 0 72352 0 -1 47040
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_638
timestamp 1669390400
transform 1 0 72800 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_55_641
timestamp 1669390400
transform 1 0 73136 0 -1 47040
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_55_673
timestamp 1669390400
transform 1 0 76720 0 -1 47040
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_55_681
timestamp 1669390400
transform 1 0 77616 0 -1 47040
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_685
timestamp 1669390400
transform 1 0 78064 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_687
timestamp 1669390400
transform 1 0 78288 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_56_2
timestamp 1669390400
transform 1 0 1568 0 1 47040
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_34
timestamp 1669390400
transform 1 0 5152 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_37
timestamp 1669390400
transform 1 0 5488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_56_101
timestamp 1669390400
transform 1 0 12656 0 1 47040
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_105
timestamp 1669390400
transform 1 0 13104 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_108
timestamp 1669390400
transform 1 0 13440 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_56_172
timestamp 1669390400
transform 1 0 20608 0 1 47040
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_176
timestamp 1669390400
transform 1 0 21056 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_179
timestamp 1669390400
transform 1 0 21392 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_56_243
timestamp 1669390400
transform 1 0 28560 0 1 47040
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_247
timestamp 1669390400
transform 1 0 29008 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_250
timestamp 1669390400
transform 1 0 29344 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_56_314
timestamp 1669390400
transform 1 0 36512 0 1 47040
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_318
timestamp 1669390400
transform 1 0 36960 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_321
timestamp 1669390400
transform 1 0 37296 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_56_385
timestamp 1669390400
transform 1 0 44464 0 1 47040
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_389
timestamp 1669390400
transform 1 0 44912 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_392
timestamp 1669390400
transform 1 0 45248 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_56_456
timestamp 1669390400
transform 1 0 52416 0 1 47040
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_460
timestamp 1669390400
transform 1 0 52864 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_463
timestamp 1669390400
transform 1 0 53200 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_56_527
timestamp 1669390400
transform 1 0 60368 0 1 47040
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_531
timestamp 1669390400
transform 1 0 60816 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_534
timestamp 1669390400
transform 1 0 61152 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_56_598
timestamp 1669390400
transform 1 0 68320 0 1 47040
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_602
timestamp 1669390400
transform 1 0 68768 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_605
timestamp 1669390400
transform 1 0 69104 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_56_669
timestamp 1669390400
transform 1 0 76272 0 1 47040
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_673
timestamp 1669390400
transform 1 0 76720 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_56_676
timestamp 1669390400
transform 1 0 77056 0 1 47040
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_56_684
timestamp 1669390400
transform 1 0 77952 0 1 47040
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_2
timestamp 1669390400
transform 1 0 1568 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_57_66
timestamp 1669390400
transform 1 0 8736 0 -1 48608
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_70
timestamp 1669390400
transform 1 0 9184 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_73
timestamp 1669390400
transform 1 0 9520 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_57_137
timestamp 1669390400
transform 1 0 16688 0 -1 48608
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_141
timestamp 1669390400
transform 1 0 17136 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_144
timestamp 1669390400
transform 1 0 17472 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_57_208
timestamp 1669390400
transform 1 0 24640 0 -1 48608
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_212
timestamp 1669390400
transform 1 0 25088 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_215
timestamp 1669390400
transform 1 0 25424 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_57_279
timestamp 1669390400
transform 1 0 32592 0 -1 48608
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_283
timestamp 1669390400
transform 1 0 33040 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_286
timestamp 1669390400
transform 1 0 33376 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_57_350
timestamp 1669390400
transform 1 0 40544 0 -1 48608
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_354
timestamp 1669390400
transform 1 0 40992 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_357
timestamp 1669390400
transform 1 0 41328 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_57_421
timestamp 1669390400
transform 1 0 48496 0 -1 48608
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_425
timestamp 1669390400
transform 1 0 48944 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_428
timestamp 1669390400
transform 1 0 49280 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_57_492
timestamp 1669390400
transform 1 0 56448 0 -1 48608
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_496
timestamp 1669390400
transform 1 0 56896 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_499
timestamp 1669390400
transform 1 0 57232 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_57_563
timestamp 1669390400
transform 1 0 64400 0 -1 48608
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_567
timestamp 1669390400
transform 1 0 64848 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_570
timestamp 1669390400
transform 1 0 65184 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_57_634
timestamp 1669390400
transform 1 0 72352 0 -1 48608
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_638
timestamp 1669390400
transform 1 0 72800 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_57_641
timestamp 1669390400
transform 1 0 73136 0 -1 48608
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_57_673
timestamp 1669390400
transform 1 0 76720 0 -1 48608
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_57_681
timestamp 1669390400
transform 1 0 77616 0 -1 48608
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_685
timestamp 1669390400
transform 1 0 78064 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_687
timestamp 1669390400
transform 1 0 78288 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_58_2
timestamp 1669390400
transform 1 0 1568 0 1 48608
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_34
timestamp 1669390400
transform 1 0 5152 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_37
timestamp 1669390400
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_58_101
timestamp 1669390400
transform 1 0 12656 0 1 48608
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_105
timestamp 1669390400
transform 1 0 13104 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_108
timestamp 1669390400
transform 1 0 13440 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_58_172
timestamp 1669390400
transform 1 0 20608 0 1 48608
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_176
timestamp 1669390400
transform 1 0 21056 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_179
timestamp 1669390400
transform 1 0 21392 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_58_243
timestamp 1669390400
transform 1 0 28560 0 1 48608
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_247
timestamp 1669390400
transform 1 0 29008 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_250
timestamp 1669390400
transform 1 0 29344 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_58_314
timestamp 1669390400
transform 1 0 36512 0 1 48608
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_318
timestamp 1669390400
transform 1 0 36960 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_321
timestamp 1669390400
transform 1 0 37296 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_58_385
timestamp 1669390400
transform 1 0 44464 0 1 48608
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_389
timestamp 1669390400
transform 1 0 44912 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_392
timestamp 1669390400
transform 1 0 45248 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_58_456
timestamp 1669390400
transform 1 0 52416 0 1 48608
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_460
timestamp 1669390400
transform 1 0 52864 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_463
timestamp 1669390400
transform 1 0 53200 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_58_527
timestamp 1669390400
transform 1 0 60368 0 1 48608
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_531
timestamp 1669390400
transform 1 0 60816 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_534
timestamp 1669390400
transform 1 0 61152 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_58_598
timestamp 1669390400
transform 1 0 68320 0 1 48608
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_602
timestamp 1669390400
transform 1 0 68768 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_605
timestamp 1669390400
transform 1 0 69104 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_58_669
timestamp 1669390400
transform 1 0 76272 0 1 48608
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_673
timestamp 1669390400
transform 1 0 76720 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_58_676
timestamp 1669390400
transform 1 0 77056 0 1 48608
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_58_684
timestamp 1669390400
transform 1 0 77952 0 1 48608
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_2
timestamp 1669390400
transform 1 0 1568 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_59_66
timestamp 1669390400
transform 1 0 8736 0 -1 50176
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_70
timestamp 1669390400
transform 1 0 9184 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_73
timestamp 1669390400
transform 1 0 9520 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_59_137
timestamp 1669390400
transform 1 0 16688 0 -1 50176
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_141
timestamp 1669390400
transform 1 0 17136 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_144
timestamp 1669390400
transform 1 0 17472 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_59_208
timestamp 1669390400
transform 1 0 24640 0 -1 50176
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_212
timestamp 1669390400
transform 1 0 25088 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_215
timestamp 1669390400
transform 1 0 25424 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_59_279
timestamp 1669390400
transform 1 0 32592 0 -1 50176
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_283
timestamp 1669390400
transform 1 0 33040 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_286
timestamp 1669390400
transform 1 0 33376 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_59_350
timestamp 1669390400
transform 1 0 40544 0 -1 50176
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_354
timestamp 1669390400
transform 1 0 40992 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_357
timestamp 1669390400
transform 1 0 41328 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_59_421
timestamp 1669390400
transform 1 0 48496 0 -1 50176
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_425
timestamp 1669390400
transform 1 0 48944 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_428
timestamp 1669390400
transform 1 0 49280 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_59_492
timestamp 1669390400
transform 1 0 56448 0 -1 50176
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_496
timestamp 1669390400
transform 1 0 56896 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_499
timestamp 1669390400
transform 1 0 57232 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_59_563
timestamp 1669390400
transform 1 0 64400 0 -1 50176
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_567
timestamp 1669390400
transform 1 0 64848 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_570
timestamp 1669390400
transform 1 0 65184 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_59_634
timestamp 1669390400
transform 1 0 72352 0 -1 50176
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_638
timestamp 1669390400
transform 1 0 72800 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_59_641
timestamp 1669390400
transform 1 0 73136 0 -1 50176
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_59_673
timestamp 1669390400
transform 1 0 76720 0 -1 50176
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_59_681
timestamp 1669390400
transform 1 0 77616 0 -1 50176
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_685
timestamp 1669390400
transform 1 0 78064 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_687
timestamp 1669390400
transform 1 0 78288 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_60_2
timestamp 1669390400
transform 1 0 1568 0 1 50176
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_34
timestamp 1669390400
transform 1 0 5152 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_37
timestamp 1669390400
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_60_101
timestamp 1669390400
transform 1 0 12656 0 1 50176
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_105
timestamp 1669390400
transform 1 0 13104 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_108
timestamp 1669390400
transform 1 0 13440 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_60_172
timestamp 1669390400
transform 1 0 20608 0 1 50176
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_176
timestamp 1669390400
transform 1 0 21056 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_179
timestamp 1669390400
transform 1 0 21392 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_60_243
timestamp 1669390400
transform 1 0 28560 0 1 50176
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_247
timestamp 1669390400
transform 1 0 29008 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_250
timestamp 1669390400
transform 1 0 29344 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_60_314
timestamp 1669390400
transform 1 0 36512 0 1 50176
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_318
timestamp 1669390400
transform 1 0 36960 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_321
timestamp 1669390400
transform 1 0 37296 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_60_385
timestamp 1669390400
transform 1 0 44464 0 1 50176
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_389
timestamp 1669390400
transform 1 0 44912 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_392
timestamp 1669390400
transform 1 0 45248 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_60_456
timestamp 1669390400
transform 1 0 52416 0 1 50176
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_460
timestamp 1669390400
transform 1 0 52864 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_463
timestamp 1669390400
transform 1 0 53200 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_60_527
timestamp 1669390400
transform 1 0 60368 0 1 50176
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_531
timestamp 1669390400
transform 1 0 60816 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_534
timestamp 1669390400
transform 1 0 61152 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_60_598
timestamp 1669390400
transform 1 0 68320 0 1 50176
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_602
timestamp 1669390400
transform 1 0 68768 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_605
timestamp 1669390400
transform 1 0 69104 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_60_669
timestamp 1669390400
transform 1 0 76272 0 1 50176
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_673
timestamp 1669390400
transform 1 0 76720 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_60_676
timestamp 1669390400
transform 1 0 77056 0 1 50176
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_60_684
timestamp 1669390400
transform 1 0 77952 0 1 50176
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_2
timestamp 1669390400
transform 1 0 1568 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_61_66
timestamp 1669390400
transform 1 0 8736 0 -1 51744
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_70
timestamp 1669390400
transform 1 0 9184 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_73
timestamp 1669390400
transform 1 0 9520 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_61_137
timestamp 1669390400
transform 1 0 16688 0 -1 51744
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_141
timestamp 1669390400
transform 1 0 17136 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_144
timestamp 1669390400
transform 1 0 17472 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_61_208
timestamp 1669390400
transform 1 0 24640 0 -1 51744
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_212
timestamp 1669390400
transform 1 0 25088 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_215
timestamp 1669390400
transform 1 0 25424 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_61_279
timestamp 1669390400
transform 1 0 32592 0 -1 51744
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_283
timestamp 1669390400
transform 1 0 33040 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_286
timestamp 1669390400
transform 1 0 33376 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_61_350
timestamp 1669390400
transform 1 0 40544 0 -1 51744
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_354
timestamp 1669390400
transform 1 0 40992 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_357
timestamp 1669390400
transform 1 0 41328 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_61_421
timestamp 1669390400
transform 1 0 48496 0 -1 51744
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_425
timestamp 1669390400
transform 1 0 48944 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_428
timestamp 1669390400
transform 1 0 49280 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_61_492
timestamp 1669390400
transform 1 0 56448 0 -1 51744
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_496
timestamp 1669390400
transform 1 0 56896 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_499
timestamp 1669390400
transform 1 0 57232 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_61_563
timestamp 1669390400
transform 1 0 64400 0 -1 51744
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_567
timestamp 1669390400
transform 1 0 64848 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_570
timestamp 1669390400
transform 1 0 65184 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_61_634
timestamp 1669390400
transform 1 0 72352 0 -1 51744
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_638
timestamp 1669390400
transform 1 0 72800 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_61_641
timestamp 1669390400
transform 1 0 73136 0 -1 51744
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_61_673
timestamp 1669390400
transform 1 0 76720 0 -1 51744
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_61_681
timestamp 1669390400
transform 1 0 77616 0 -1 51744
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_685
timestamp 1669390400
transform 1 0 78064 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_687
timestamp 1669390400
transform 1 0 78288 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_62_2
timestamp 1669390400
transform 1 0 1568 0 1 51744
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_34
timestamp 1669390400
transform 1 0 5152 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_37
timestamp 1669390400
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_62_101
timestamp 1669390400
transform 1 0 12656 0 1 51744
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_105
timestamp 1669390400
transform 1 0 13104 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_108
timestamp 1669390400
transform 1 0 13440 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_62_172
timestamp 1669390400
transform 1 0 20608 0 1 51744
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_176
timestamp 1669390400
transform 1 0 21056 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_179
timestamp 1669390400
transform 1 0 21392 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_62_243
timestamp 1669390400
transform 1 0 28560 0 1 51744
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_247
timestamp 1669390400
transform 1 0 29008 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_250
timestamp 1669390400
transform 1 0 29344 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_62_314
timestamp 1669390400
transform 1 0 36512 0 1 51744
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_318
timestamp 1669390400
transform 1 0 36960 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_321
timestamp 1669390400
transform 1 0 37296 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_62_385
timestamp 1669390400
transform 1 0 44464 0 1 51744
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_389
timestamp 1669390400
transform 1 0 44912 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_392
timestamp 1669390400
transform 1 0 45248 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_62_456
timestamp 1669390400
transform 1 0 52416 0 1 51744
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_460
timestamp 1669390400
transform 1 0 52864 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_463
timestamp 1669390400
transform 1 0 53200 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_62_527
timestamp 1669390400
transform 1 0 60368 0 1 51744
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_531
timestamp 1669390400
transform 1 0 60816 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_534
timestamp 1669390400
transform 1 0 61152 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_62_598
timestamp 1669390400
transform 1 0 68320 0 1 51744
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_602
timestamp 1669390400
transform 1 0 68768 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_605
timestamp 1669390400
transform 1 0 69104 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_62_669
timestamp 1669390400
transform 1 0 76272 0 1 51744
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_673
timestamp 1669390400
transform 1 0 76720 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_62_676
timestamp 1669390400
transform 1 0 77056 0 1 51744
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_62_684
timestamp 1669390400
transform 1 0 77952 0 1 51744
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_2
timestamp 1669390400
transform 1 0 1568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_63_66
timestamp 1669390400
transform 1 0 8736 0 -1 53312
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_70
timestamp 1669390400
transform 1 0 9184 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_73
timestamp 1669390400
transform 1 0 9520 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_63_137
timestamp 1669390400
transform 1 0 16688 0 -1 53312
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_141
timestamp 1669390400
transform 1 0 17136 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_144
timestamp 1669390400
transform 1 0 17472 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_63_208
timestamp 1669390400
transform 1 0 24640 0 -1 53312
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_212
timestamp 1669390400
transform 1 0 25088 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_215
timestamp 1669390400
transform 1 0 25424 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_63_279
timestamp 1669390400
transform 1 0 32592 0 -1 53312
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_283
timestamp 1669390400
transform 1 0 33040 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_286
timestamp 1669390400
transform 1 0 33376 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_63_350
timestamp 1669390400
transform 1 0 40544 0 -1 53312
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_354
timestamp 1669390400
transform 1 0 40992 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_357
timestamp 1669390400
transform 1 0 41328 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_63_421
timestamp 1669390400
transform 1 0 48496 0 -1 53312
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_425
timestamp 1669390400
transform 1 0 48944 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_428
timestamp 1669390400
transform 1 0 49280 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_63_492
timestamp 1669390400
transform 1 0 56448 0 -1 53312
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_496
timestamp 1669390400
transform 1 0 56896 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_499
timestamp 1669390400
transform 1 0 57232 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_63_563
timestamp 1669390400
transform 1 0 64400 0 -1 53312
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_567
timestamp 1669390400
transform 1 0 64848 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_570
timestamp 1669390400
transform 1 0 65184 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_63_634
timestamp 1669390400
transform 1 0 72352 0 -1 53312
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_638
timestamp 1669390400
transform 1 0 72800 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_63_641
timestamp 1669390400
transform 1 0 73136 0 -1 53312
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_63_673
timestamp 1669390400
transform 1 0 76720 0 -1 53312
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_63_681
timestamp 1669390400
transform 1 0 77616 0 -1 53312
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_685
timestamp 1669390400
transform 1 0 78064 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_687
timestamp 1669390400
transform 1 0 78288 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_64_2
timestamp 1669390400
transform 1 0 1568 0 1 53312
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_34
timestamp 1669390400
transform 1 0 5152 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_37
timestamp 1669390400
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_64_101
timestamp 1669390400
transform 1 0 12656 0 1 53312
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_105
timestamp 1669390400
transform 1 0 13104 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_108
timestamp 1669390400
transform 1 0 13440 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_64_172
timestamp 1669390400
transform 1 0 20608 0 1 53312
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_176
timestamp 1669390400
transform 1 0 21056 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_179
timestamp 1669390400
transform 1 0 21392 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_64_243
timestamp 1669390400
transform 1 0 28560 0 1 53312
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_247
timestamp 1669390400
transform 1 0 29008 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_250
timestamp 1669390400
transform 1 0 29344 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_64_314
timestamp 1669390400
transform 1 0 36512 0 1 53312
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_318
timestamp 1669390400
transform 1 0 36960 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_321
timestamp 1669390400
transform 1 0 37296 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_64_385
timestamp 1669390400
transform 1 0 44464 0 1 53312
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_389
timestamp 1669390400
transform 1 0 44912 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_392
timestamp 1669390400
transform 1 0 45248 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_64_456
timestamp 1669390400
transform 1 0 52416 0 1 53312
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_460
timestamp 1669390400
transform 1 0 52864 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_463
timestamp 1669390400
transform 1 0 53200 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_64_527
timestamp 1669390400
transform 1 0 60368 0 1 53312
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_531
timestamp 1669390400
transform 1 0 60816 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_534
timestamp 1669390400
transform 1 0 61152 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_64_598
timestamp 1669390400
transform 1 0 68320 0 1 53312
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_602
timestamp 1669390400
transform 1 0 68768 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_605
timestamp 1669390400
transform 1 0 69104 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_64_669
timestamp 1669390400
transform 1 0 76272 0 1 53312
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_673
timestamp 1669390400
transform 1 0 76720 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_64_676
timestamp 1669390400
transform 1 0 77056 0 1 53312
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_64_684
timestamp 1669390400
transform 1 0 77952 0 1 53312
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_2
timestamp 1669390400
transform 1 0 1568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_65_66
timestamp 1669390400
transform 1 0 8736 0 -1 54880
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_70
timestamp 1669390400
transform 1 0 9184 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_73
timestamp 1669390400
transform 1 0 9520 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_65_137
timestamp 1669390400
transform 1 0 16688 0 -1 54880
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_141
timestamp 1669390400
transform 1 0 17136 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_144
timestamp 1669390400
transform 1 0 17472 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_65_208
timestamp 1669390400
transform 1 0 24640 0 -1 54880
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_212
timestamp 1669390400
transform 1 0 25088 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_215
timestamp 1669390400
transform 1 0 25424 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_65_279
timestamp 1669390400
transform 1 0 32592 0 -1 54880
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_283
timestamp 1669390400
transform 1 0 33040 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_286
timestamp 1669390400
transform 1 0 33376 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_65_350
timestamp 1669390400
transform 1 0 40544 0 -1 54880
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_354
timestamp 1669390400
transform 1 0 40992 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_357
timestamp 1669390400
transform 1 0 41328 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_65_421
timestamp 1669390400
transform 1 0 48496 0 -1 54880
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_425
timestamp 1669390400
transform 1 0 48944 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_428
timestamp 1669390400
transform 1 0 49280 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_65_492
timestamp 1669390400
transform 1 0 56448 0 -1 54880
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_496
timestamp 1669390400
transform 1 0 56896 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_499
timestamp 1669390400
transform 1 0 57232 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_65_563
timestamp 1669390400
transform 1 0 64400 0 -1 54880
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_567
timestamp 1669390400
transform 1 0 64848 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_570
timestamp 1669390400
transform 1 0 65184 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_65_634
timestamp 1669390400
transform 1 0 72352 0 -1 54880
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_638
timestamp 1669390400
transform 1 0 72800 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_65_641
timestamp 1669390400
transform 1 0 73136 0 -1 54880
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_65_673
timestamp 1669390400
transform 1 0 76720 0 -1 54880
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_65_681
timestamp 1669390400
transform 1 0 77616 0 -1 54880
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_685
timestamp 1669390400
transform 1 0 78064 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_687
timestamp 1669390400
transform 1 0 78288 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_66_2
timestamp 1669390400
transform 1 0 1568 0 1 54880
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_34
timestamp 1669390400
transform 1 0 5152 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_37
timestamp 1669390400
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_66_101
timestamp 1669390400
transform 1 0 12656 0 1 54880
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_105
timestamp 1669390400
transform 1 0 13104 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_108
timestamp 1669390400
transform 1 0 13440 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_66_172
timestamp 1669390400
transform 1 0 20608 0 1 54880
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_176
timestamp 1669390400
transform 1 0 21056 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_179
timestamp 1669390400
transform 1 0 21392 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_66_243
timestamp 1669390400
transform 1 0 28560 0 1 54880
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_247
timestamp 1669390400
transform 1 0 29008 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_250
timestamp 1669390400
transform 1 0 29344 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_66_314
timestamp 1669390400
transform 1 0 36512 0 1 54880
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_318
timestamp 1669390400
transform 1 0 36960 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_321
timestamp 1669390400
transform 1 0 37296 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_66_385
timestamp 1669390400
transform 1 0 44464 0 1 54880
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_389
timestamp 1669390400
transform 1 0 44912 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_392
timestamp 1669390400
transform 1 0 45248 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_66_456
timestamp 1669390400
transform 1 0 52416 0 1 54880
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_460
timestamp 1669390400
transform 1 0 52864 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_463
timestamp 1669390400
transform 1 0 53200 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_66_527
timestamp 1669390400
transform 1 0 60368 0 1 54880
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_531
timestamp 1669390400
transform 1 0 60816 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_534
timestamp 1669390400
transform 1 0 61152 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_66_598
timestamp 1669390400
transform 1 0 68320 0 1 54880
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_602
timestamp 1669390400
transform 1 0 68768 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_605
timestamp 1669390400
transform 1 0 69104 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_66_669
timestamp 1669390400
transform 1 0 76272 0 1 54880
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_673
timestamp 1669390400
transform 1 0 76720 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_66_676
timestamp 1669390400
transform 1 0 77056 0 1 54880
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_66_684
timestamp 1669390400
transform 1 0 77952 0 1 54880
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_2
timestamp 1669390400
transform 1 0 1568 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_67_66
timestamp 1669390400
transform 1 0 8736 0 -1 56448
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_70
timestamp 1669390400
transform 1 0 9184 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_73
timestamp 1669390400
transform 1 0 9520 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_67_137
timestamp 1669390400
transform 1 0 16688 0 -1 56448
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_141
timestamp 1669390400
transform 1 0 17136 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_144
timestamp 1669390400
transform 1 0 17472 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_67_208
timestamp 1669390400
transform 1 0 24640 0 -1 56448
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_212
timestamp 1669390400
transform 1 0 25088 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_215
timestamp 1669390400
transform 1 0 25424 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_67_279
timestamp 1669390400
transform 1 0 32592 0 -1 56448
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_283
timestamp 1669390400
transform 1 0 33040 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_286
timestamp 1669390400
transform 1 0 33376 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_67_350
timestamp 1669390400
transform 1 0 40544 0 -1 56448
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_354
timestamp 1669390400
transform 1 0 40992 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_357
timestamp 1669390400
transform 1 0 41328 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_67_421
timestamp 1669390400
transform 1 0 48496 0 -1 56448
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_425
timestamp 1669390400
transform 1 0 48944 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_428
timestamp 1669390400
transform 1 0 49280 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_67_492
timestamp 1669390400
transform 1 0 56448 0 -1 56448
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_496
timestamp 1669390400
transform 1 0 56896 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_499
timestamp 1669390400
transform 1 0 57232 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_67_563
timestamp 1669390400
transform 1 0 64400 0 -1 56448
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_567
timestamp 1669390400
transform 1 0 64848 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_570
timestamp 1669390400
transform 1 0 65184 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_67_634
timestamp 1669390400
transform 1 0 72352 0 -1 56448
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_638
timestamp 1669390400
transform 1 0 72800 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_67_641
timestamp 1669390400
transform 1 0 73136 0 -1 56448
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_67_673
timestamp 1669390400
transform 1 0 76720 0 -1 56448
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_67_681
timestamp 1669390400
transform 1 0 77616 0 -1 56448
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_685
timestamp 1669390400
transform 1 0 78064 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_687
timestamp 1669390400
transform 1 0 78288 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_68_2
timestamp 1669390400
transform 1 0 1568 0 1 56448
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_34
timestamp 1669390400
transform 1 0 5152 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_37
timestamp 1669390400
transform 1 0 5488 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_68_101
timestamp 1669390400
transform 1 0 12656 0 1 56448
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_105
timestamp 1669390400
transform 1 0 13104 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_108
timestamp 1669390400
transform 1 0 13440 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_68_172
timestamp 1669390400
transform 1 0 20608 0 1 56448
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_176
timestamp 1669390400
transform 1 0 21056 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_179
timestamp 1669390400
transform 1 0 21392 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_68_243
timestamp 1669390400
transform 1 0 28560 0 1 56448
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_247
timestamp 1669390400
transform 1 0 29008 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_250
timestamp 1669390400
transform 1 0 29344 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_68_314
timestamp 1669390400
transform 1 0 36512 0 1 56448
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_318
timestamp 1669390400
transform 1 0 36960 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_321
timestamp 1669390400
transform 1 0 37296 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_68_385
timestamp 1669390400
transform 1 0 44464 0 1 56448
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_389
timestamp 1669390400
transform 1 0 44912 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_392
timestamp 1669390400
transform 1 0 45248 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_68_456
timestamp 1669390400
transform 1 0 52416 0 1 56448
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_460
timestamp 1669390400
transform 1 0 52864 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_463
timestamp 1669390400
transform 1 0 53200 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_68_527
timestamp 1669390400
transform 1 0 60368 0 1 56448
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_531
timestamp 1669390400
transform 1 0 60816 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_534
timestamp 1669390400
transform 1 0 61152 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_68_598
timestamp 1669390400
transform 1 0 68320 0 1 56448
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_602
timestamp 1669390400
transform 1 0 68768 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_605
timestamp 1669390400
transform 1 0 69104 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_68_669
timestamp 1669390400
transform 1 0 76272 0 1 56448
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_673
timestamp 1669390400
transform 1 0 76720 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_68_676
timestamp 1669390400
transform 1 0 77056 0 1 56448
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_68_684
timestamp 1669390400
transform 1 0 77952 0 1 56448
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_2
timestamp 1669390400
transform 1 0 1568 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_69_66
timestamp 1669390400
transform 1 0 8736 0 -1 58016
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_70
timestamp 1669390400
transform 1 0 9184 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_73
timestamp 1669390400
transform 1 0 9520 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_69_137
timestamp 1669390400
transform 1 0 16688 0 -1 58016
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_141
timestamp 1669390400
transform 1 0 17136 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_144
timestamp 1669390400
transform 1 0 17472 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_69_208
timestamp 1669390400
transform 1 0 24640 0 -1 58016
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_212
timestamp 1669390400
transform 1 0 25088 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_215
timestamp 1669390400
transform 1 0 25424 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_69_279
timestamp 1669390400
transform 1 0 32592 0 -1 58016
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_283
timestamp 1669390400
transform 1 0 33040 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_286
timestamp 1669390400
transform 1 0 33376 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_69_350
timestamp 1669390400
transform 1 0 40544 0 -1 58016
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_354
timestamp 1669390400
transform 1 0 40992 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_357
timestamp 1669390400
transform 1 0 41328 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_69_421
timestamp 1669390400
transform 1 0 48496 0 -1 58016
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_425
timestamp 1669390400
transform 1 0 48944 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_428
timestamp 1669390400
transform 1 0 49280 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_69_492
timestamp 1669390400
transform 1 0 56448 0 -1 58016
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_496
timestamp 1669390400
transform 1 0 56896 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_499
timestamp 1669390400
transform 1 0 57232 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_69_563
timestamp 1669390400
transform 1 0 64400 0 -1 58016
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_567
timestamp 1669390400
transform 1 0 64848 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_570
timestamp 1669390400
transform 1 0 65184 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_69_634
timestamp 1669390400
transform 1 0 72352 0 -1 58016
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_638
timestamp 1669390400
transform 1 0 72800 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_69_641
timestamp 1669390400
transform 1 0 73136 0 -1 58016
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_69_673
timestamp 1669390400
transform 1 0 76720 0 -1 58016
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_69_681
timestamp 1669390400
transform 1 0 77616 0 -1 58016
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_685
timestamp 1669390400
transform 1 0 78064 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_687
timestamp 1669390400
transform 1 0 78288 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_70_2
timestamp 1669390400
transform 1 0 1568 0 1 58016
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_34
timestamp 1669390400
transform 1 0 5152 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_37
timestamp 1669390400
transform 1 0 5488 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_70_101
timestamp 1669390400
transform 1 0 12656 0 1 58016
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_105
timestamp 1669390400
transform 1 0 13104 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_108
timestamp 1669390400
transform 1 0 13440 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_70_172
timestamp 1669390400
transform 1 0 20608 0 1 58016
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_176
timestamp 1669390400
transform 1 0 21056 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_179
timestamp 1669390400
transform 1 0 21392 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_70_243
timestamp 1669390400
transform 1 0 28560 0 1 58016
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_247
timestamp 1669390400
transform 1 0 29008 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_250
timestamp 1669390400
transform 1 0 29344 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_70_314
timestamp 1669390400
transform 1 0 36512 0 1 58016
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_318
timestamp 1669390400
transform 1 0 36960 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_321
timestamp 1669390400
transform 1 0 37296 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_70_385
timestamp 1669390400
transform 1 0 44464 0 1 58016
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_389
timestamp 1669390400
transform 1 0 44912 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_392
timestamp 1669390400
transform 1 0 45248 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_70_456
timestamp 1669390400
transform 1 0 52416 0 1 58016
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_460
timestamp 1669390400
transform 1 0 52864 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_463
timestamp 1669390400
transform 1 0 53200 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_70_527
timestamp 1669390400
transform 1 0 60368 0 1 58016
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_531
timestamp 1669390400
transform 1 0 60816 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_534
timestamp 1669390400
transform 1 0 61152 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_70_598
timestamp 1669390400
transform 1 0 68320 0 1 58016
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_602
timestamp 1669390400
transform 1 0 68768 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_605
timestamp 1669390400
transform 1 0 69104 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_70_669
timestamp 1669390400
transform 1 0 76272 0 1 58016
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_673
timestamp 1669390400
transform 1 0 76720 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_70_676
timestamp 1669390400
transform 1 0 77056 0 1 58016
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_70_684
timestamp 1669390400
transform 1 0 77952 0 1 58016
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_2
timestamp 1669390400
transform 1 0 1568 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_71_66
timestamp 1669390400
transform 1 0 8736 0 -1 59584
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_70
timestamp 1669390400
transform 1 0 9184 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_73
timestamp 1669390400
transform 1 0 9520 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_71_137
timestamp 1669390400
transform 1 0 16688 0 -1 59584
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_141
timestamp 1669390400
transform 1 0 17136 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_144
timestamp 1669390400
transform 1 0 17472 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_71_208
timestamp 1669390400
transform 1 0 24640 0 -1 59584
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_212
timestamp 1669390400
transform 1 0 25088 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_215
timestamp 1669390400
transform 1 0 25424 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_71_279
timestamp 1669390400
transform 1 0 32592 0 -1 59584
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_283
timestamp 1669390400
transform 1 0 33040 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_286
timestamp 1669390400
transform 1 0 33376 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_71_350
timestamp 1669390400
transform 1 0 40544 0 -1 59584
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_354
timestamp 1669390400
transform 1 0 40992 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_357
timestamp 1669390400
transform 1 0 41328 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_71_421
timestamp 1669390400
transform 1 0 48496 0 -1 59584
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_425
timestamp 1669390400
transform 1 0 48944 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_428
timestamp 1669390400
transform 1 0 49280 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_71_492
timestamp 1669390400
transform 1 0 56448 0 -1 59584
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_496
timestamp 1669390400
transform 1 0 56896 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_499
timestamp 1669390400
transform 1 0 57232 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_71_563
timestamp 1669390400
transform 1 0 64400 0 -1 59584
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_567
timestamp 1669390400
transform 1 0 64848 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_570
timestamp 1669390400
transform 1 0 65184 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_71_634
timestamp 1669390400
transform 1 0 72352 0 -1 59584
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_638
timestamp 1669390400
transform 1 0 72800 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_71_641
timestamp 1669390400
transform 1 0 73136 0 -1 59584
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_71_673
timestamp 1669390400
transform 1 0 76720 0 -1 59584
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_71_681
timestamp 1669390400
transform 1 0 77616 0 -1 59584
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_685
timestamp 1669390400
transform 1 0 78064 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_687
timestamp 1669390400
transform 1 0 78288 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_72_2
timestamp 1669390400
transform 1 0 1568 0 1 59584
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_34
timestamp 1669390400
transform 1 0 5152 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_37
timestamp 1669390400
transform 1 0 5488 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_72_101
timestamp 1669390400
transform 1 0 12656 0 1 59584
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_105
timestamp 1669390400
transform 1 0 13104 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_108
timestamp 1669390400
transform 1 0 13440 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_72_172
timestamp 1669390400
transform 1 0 20608 0 1 59584
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_176
timestamp 1669390400
transform 1 0 21056 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_179
timestamp 1669390400
transform 1 0 21392 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_72_243
timestamp 1669390400
transform 1 0 28560 0 1 59584
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_247
timestamp 1669390400
transform 1 0 29008 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_250
timestamp 1669390400
transform 1 0 29344 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_72_314
timestamp 1669390400
transform 1 0 36512 0 1 59584
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_318
timestamp 1669390400
transform 1 0 36960 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_321
timestamp 1669390400
transform 1 0 37296 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_72_385
timestamp 1669390400
transform 1 0 44464 0 1 59584
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_389
timestamp 1669390400
transform 1 0 44912 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_392
timestamp 1669390400
transform 1 0 45248 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_72_456
timestamp 1669390400
transform 1 0 52416 0 1 59584
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_460
timestamp 1669390400
transform 1 0 52864 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_463
timestamp 1669390400
transform 1 0 53200 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_72_527
timestamp 1669390400
transform 1 0 60368 0 1 59584
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_531
timestamp 1669390400
transform 1 0 60816 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_534
timestamp 1669390400
transform 1 0 61152 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_72_598
timestamp 1669390400
transform 1 0 68320 0 1 59584
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_602
timestamp 1669390400
transform 1 0 68768 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_605
timestamp 1669390400
transform 1 0 69104 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_72_669
timestamp 1669390400
transform 1 0 76272 0 1 59584
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_673
timestamp 1669390400
transform 1 0 76720 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_72_676
timestamp 1669390400
transform 1 0 77056 0 1 59584
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_72_684
timestamp 1669390400
transform 1 0 77952 0 1 59584
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_2
timestamp 1669390400
transform 1 0 1568 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_73_66
timestamp 1669390400
transform 1 0 8736 0 -1 61152
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_70
timestamp 1669390400
transform 1 0 9184 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_73
timestamp 1669390400
transform 1 0 9520 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_73_137
timestamp 1669390400
transform 1 0 16688 0 -1 61152
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_141
timestamp 1669390400
transform 1 0 17136 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_144
timestamp 1669390400
transform 1 0 17472 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_73_208
timestamp 1669390400
transform 1 0 24640 0 -1 61152
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_212
timestamp 1669390400
transform 1 0 25088 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_215
timestamp 1669390400
transform 1 0 25424 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_73_279
timestamp 1669390400
transform 1 0 32592 0 -1 61152
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_283
timestamp 1669390400
transform 1 0 33040 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_286
timestamp 1669390400
transform 1 0 33376 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_73_350
timestamp 1669390400
transform 1 0 40544 0 -1 61152
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_354
timestamp 1669390400
transform 1 0 40992 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_357
timestamp 1669390400
transform 1 0 41328 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_73_421
timestamp 1669390400
transform 1 0 48496 0 -1 61152
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_425
timestamp 1669390400
transform 1 0 48944 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_428
timestamp 1669390400
transform 1 0 49280 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_73_492
timestamp 1669390400
transform 1 0 56448 0 -1 61152
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_496
timestamp 1669390400
transform 1 0 56896 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_499
timestamp 1669390400
transform 1 0 57232 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_73_563
timestamp 1669390400
transform 1 0 64400 0 -1 61152
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_567
timestamp 1669390400
transform 1 0 64848 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_570
timestamp 1669390400
transform 1 0 65184 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_73_634
timestamp 1669390400
transform 1 0 72352 0 -1 61152
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_638
timestamp 1669390400
transform 1 0 72800 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_73_641
timestamp 1669390400
transform 1 0 73136 0 -1 61152
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_73_673
timestamp 1669390400
transform 1 0 76720 0 -1 61152
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_73_681
timestamp 1669390400
transform 1 0 77616 0 -1 61152
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_685
timestamp 1669390400
transform 1 0 78064 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_687
timestamp 1669390400
transform 1 0 78288 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_74_2
timestamp 1669390400
transform 1 0 1568 0 1 61152
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_34
timestamp 1669390400
transform 1 0 5152 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_37
timestamp 1669390400
transform 1 0 5488 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_74_101
timestamp 1669390400
transform 1 0 12656 0 1 61152
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_105
timestamp 1669390400
transform 1 0 13104 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_108
timestamp 1669390400
transform 1 0 13440 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_74_172
timestamp 1669390400
transform 1 0 20608 0 1 61152
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_176
timestamp 1669390400
transform 1 0 21056 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_179
timestamp 1669390400
transform 1 0 21392 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_74_243
timestamp 1669390400
transform 1 0 28560 0 1 61152
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_247
timestamp 1669390400
transform 1 0 29008 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_250
timestamp 1669390400
transform 1 0 29344 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_74_314
timestamp 1669390400
transform 1 0 36512 0 1 61152
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_318
timestamp 1669390400
transform 1 0 36960 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_321
timestamp 1669390400
transform 1 0 37296 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_74_385
timestamp 1669390400
transform 1 0 44464 0 1 61152
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_389
timestamp 1669390400
transform 1 0 44912 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_392
timestamp 1669390400
transform 1 0 45248 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_74_456
timestamp 1669390400
transform 1 0 52416 0 1 61152
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_460
timestamp 1669390400
transform 1 0 52864 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_463
timestamp 1669390400
transform 1 0 53200 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_74_527
timestamp 1669390400
transform 1 0 60368 0 1 61152
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_531
timestamp 1669390400
transform 1 0 60816 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_534
timestamp 1669390400
transform 1 0 61152 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_74_598
timestamp 1669390400
transform 1 0 68320 0 1 61152
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_602
timestamp 1669390400
transform 1 0 68768 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_605
timestamp 1669390400
transform 1 0 69104 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_74_669
timestamp 1669390400
transform 1 0 76272 0 1 61152
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_673
timestamp 1669390400
transform 1 0 76720 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_74_676
timestamp 1669390400
transform 1 0 77056 0 1 61152
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_74_684
timestamp 1669390400
transform 1 0 77952 0 1 61152
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_2
timestamp 1669390400
transform 1 0 1568 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_75_66
timestamp 1669390400
transform 1 0 8736 0 -1 62720
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_70
timestamp 1669390400
transform 1 0 9184 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_73
timestamp 1669390400
transform 1 0 9520 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_75_137
timestamp 1669390400
transform 1 0 16688 0 -1 62720
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_141
timestamp 1669390400
transform 1 0 17136 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_144
timestamp 1669390400
transform 1 0 17472 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_75_208
timestamp 1669390400
transform 1 0 24640 0 -1 62720
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_212
timestamp 1669390400
transform 1 0 25088 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_215
timestamp 1669390400
transform 1 0 25424 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_75_279
timestamp 1669390400
transform 1 0 32592 0 -1 62720
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_283
timestamp 1669390400
transform 1 0 33040 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_286
timestamp 1669390400
transform 1 0 33376 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_75_350
timestamp 1669390400
transform 1 0 40544 0 -1 62720
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_354
timestamp 1669390400
transform 1 0 40992 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_357
timestamp 1669390400
transform 1 0 41328 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_75_421
timestamp 1669390400
transform 1 0 48496 0 -1 62720
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_425
timestamp 1669390400
transform 1 0 48944 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_428
timestamp 1669390400
transform 1 0 49280 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_75_492
timestamp 1669390400
transform 1 0 56448 0 -1 62720
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_496
timestamp 1669390400
transform 1 0 56896 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_499
timestamp 1669390400
transform 1 0 57232 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_75_563
timestamp 1669390400
transform 1 0 64400 0 -1 62720
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_567
timestamp 1669390400
transform 1 0 64848 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_570
timestamp 1669390400
transform 1 0 65184 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_75_634
timestamp 1669390400
transform 1 0 72352 0 -1 62720
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_638
timestamp 1669390400
transform 1 0 72800 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_75_641
timestamp 1669390400
transform 1 0 73136 0 -1 62720
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_75_673
timestamp 1669390400
transform 1 0 76720 0 -1 62720
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_75_681
timestamp 1669390400
transform 1 0 77616 0 -1 62720
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_685
timestamp 1669390400
transform 1 0 78064 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_687
timestamp 1669390400
transform 1 0 78288 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_76_2
timestamp 1669390400
transform 1 0 1568 0 1 62720
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_34
timestamp 1669390400
transform 1 0 5152 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_37
timestamp 1669390400
transform 1 0 5488 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_76_101
timestamp 1669390400
transform 1 0 12656 0 1 62720
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_105
timestamp 1669390400
transform 1 0 13104 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_108
timestamp 1669390400
transform 1 0 13440 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_76_172
timestamp 1669390400
transform 1 0 20608 0 1 62720
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_176
timestamp 1669390400
transform 1 0 21056 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_179
timestamp 1669390400
transform 1 0 21392 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_76_243
timestamp 1669390400
transform 1 0 28560 0 1 62720
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_247
timestamp 1669390400
transform 1 0 29008 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_250
timestamp 1669390400
transform 1 0 29344 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_76_314
timestamp 1669390400
transform 1 0 36512 0 1 62720
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_318
timestamp 1669390400
transform 1 0 36960 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_321
timestamp 1669390400
transform 1 0 37296 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_76_385
timestamp 1669390400
transform 1 0 44464 0 1 62720
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_389
timestamp 1669390400
transform 1 0 44912 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_392
timestamp 1669390400
transform 1 0 45248 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_76_456
timestamp 1669390400
transform 1 0 52416 0 1 62720
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_460
timestamp 1669390400
transform 1 0 52864 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_463
timestamp 1669390400
transform 1 0 53200 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_76_527
timestamp 1669390400
transform 1 0 60368 0 1 62720
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_531
timestamp 1669390400
transform 1 0 60816 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_534
timestamp 1669390400
transform 1 0 61152 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_76_598
timestamp 1669390400
transform 1 0 68320 0 1 62720
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_602
timestamp 1669390400
transform 1 0 68768 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_605
timestamp 1669390400
transform 1 0 69104 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_76_669
timestamp 1669390400
transform 1 0 76272 0 1 62720
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_673
timestamp 1669390400
transform 1 0 76720 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_76_676
timestamp 1669390400
transform 1 0 77056 0 1 62720
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_76_684
timestamp 1669390400
transform 1 0 77952 0 1 62720
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_2
timestamp 1669390400
transform 1 0 1568 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_77_66
timestamp 1669390400
transform 1 0 8736 0 -1 64288
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_70
timestamp 1669390400
transform 1 0 9184 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_73
timestamp 1669390400
transform 1 0 9520 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_77_137
timestamp 1669390400
transform 1 0 16688 0 -1 64288
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_141
timestamp 1669390400
transform 1 0 17136 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_144
timestamp 1669390400
transform 1 0 17472 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_77_208
timestamp 1669390400
transform 1 0 24640 0 -1 64288
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_212
timestamp 1669390400
transform 1 0 25088 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_215
timestamp 1669390400
transform 1 0 25424 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_77_279
timestamp 1669390400
transform 1 0 32592 0 -1 64288
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_283
timestamp 1669390400
transform 1 0 33040 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_286
timestamp 1669390400
transform 1 0 33376 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_77_350
timestamp 1669390400
transform 1 0 40544 0 -1 64288
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_354
timestamp 1669390400
transform 1 0 40992 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_357
timestamp 1669390400
transform 1 0 41328 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_77_421
timestamp 1669390400
transform 1 0 48496 0 -1 64288
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_425
timestamp 1669390400
transform 1 0 48944 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_428
timestamp 1669390400
transform 1 0 49280 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_77_492
timestamp 1669390400
transform 1 0 56448 0 -1 64288
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_496
timestamp 1669390400
transform 1 0 56896 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_499
timestamp 1669390400
transform 1 0 57232 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_77_563
timestamp 1669390400
transform 1 0 64400 0 -1 64288
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_567
timestamp 1669390400
transform 1 0 64848 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_570
timestamp 1669390400
transform 1 0 65184 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_77_634
timestamp 1669390400
transform 1 0 72352 0 -1 64288
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_638
timestamp 1669390400
transform 1 0 72800 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_77_641
timestamp 1669390400
transform 1 0 73136 0 -1 64288
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_77_673
timestamp 1669390400
transform 1 0 76720 0 -1 64288
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_77_681
timestamp 1669390400
transform 1 0 77616 0 -1 64288
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_685
timestamp 1669390400
transform 1 0 78064 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_687
timestamp 1669390400
transform 1 0 78288 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_78_2
timestamp 1669390400
transform 1 0 1568 0 1 64288
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_34
timestamp 1669390400
transform 1 0 5152 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_37
timestamp 1669390400
transform 1 0 5488 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_78_101
timestamp 1669390400
transform 1 0 12656 0 1 64288
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_105
timestamp 1669390400
transform 1 0 13104 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_108
timestamp 1669390400
transform 1 0 13440 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_78_172
timestamp 1669390400
transform 1 0 20608 0 1 64288
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_176
timestamp 1669390400
transform 1 0 21056 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_179
timestamp 1669390400
transform 1 0 21392 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_78_243
timestamp 1669390400
transform 1 0 28560 0 1 64288
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_247
timestamp 1669390400
transform 1 0 29008 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_250
timestamp 1669390400
transform 1 0 29344 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_78_314
timestamp 1669390400
transform 1 0 36512 0 1 64288
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_318
timestamp 1669390400
transform 1 0 36960 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_321
timestamp 1669390400
transform 1 0 37296 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_78_385
timestamp 1669390400
transform 1 0 44464 0 1 64288
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_389
timestamp 1669390400
transform 1 0 44912 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_392
timestamp 1669390400
transform 1 0 45248 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_78_456
timestamp 1669390400
transform 1 0 52416 0 1 64288
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_460
timestamp 1669390400
transform 1 0 52864 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_463
timestamp 1669390400
transform 1 0 53200 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_78_527
timestamp 1669390400
transform 1 0 60368 0 1 64288
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_531
timestamp 1669390400
transform 1 0 60816 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_534
timestamp 1669390400
transform 1 0 61152 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_78_598
timestamp 1669390400
transform 1 0 68320 0 1 64288
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_602
timestamp 1669390400
transform 1 0 68768 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_605
timestamp 1669390400
transform 1 0 69104 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_78_669
timestamp 1669390400
transform 1 0 76272 0 1 64288
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_673
timestamp 1669390400
transform 1 0 76720 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_78_676
timestamp 1669390400
transform 1 0 77056 0 1 64288
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_78_684
timestamp 1669390400
transform 1 0 77952 0 1 64288
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_2
timestamp 1669390400
transform 1 0 1568 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_79_66
timestamp 1669390400
transform 1 0 8736 0 -1 65856
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_70
timestamp 1669390400
transform 1 0 9184 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_73
timestamp 1669390400
transform 1 0 9520 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_79_137
timestamp 1669390400
transform 1 0 16688 0 -1 65856
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_141
timestamp 1669390400
transform 1 0 17136 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_144
timestamp 1669390400
transform 1 0 17472 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_79_208
timestamp 1669390400
transform 1 0 24640 0 -1 65856
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_212
timestamp 1669390400
transform 1 0 25088 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_215
timestamp 1669390400
transform 1 0 25424 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_79_279
timestamp 1669390400
transform 1 0 32592 0 -1 65856
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_283
timestamp 1669390400
transform 1 0 33040 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_286
timestamp 1669390400
transform 1 0 33376 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_79_350
timestamp 1669390400
transform 1 0 40544 0 -1 65856
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_354
timestamp 1669390400
transform 1 0 40992 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_357
timestamp 1669390400
transform 1 0 41328 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_79_421
timestamp 1669390400
transform 1 0 48496 0 -1 65856
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_425
timestamp 1669390400
transform 1 0 48944 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_428
timestamp 1669390400
transform 1 0 49280 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_79_492
timestamp 1669390400
transform 1 0 56448 0 -1 65856
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_496
timestamp 1669390400
transform 1 0 56896 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_499
timestamp 1669390400
transform 1 0 57232 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_79_563
timestamp 1669390400
transform 1 0 64400 0 -1 65856
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_567
timestamp 1669390400
transform 1 0 64848 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_570
timestamp 1669390400
transform 1 0 65184 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_79_634
timestamp 1669390400
transform 1 0 72352 0 -1 65856
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_638
timestamp 1669390400
transform 1 0 72800 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_79_641
timestamp 1669390400
transform 1 0 73136 0 -1 65856
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_79_673
timestamp 1669390400
transform 1 0 76720 0 -1 65856
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_79_681
timestamp 1669390400
transform 1 0 77616 0 -1 65856
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_685
timestamp 1669390400
transform 1 0 78064 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_687
timestamp 1669390400
transform 1 0 78288 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_80_2
timestamp 1669390400
transform 1 0 1568 0 1 65856
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_34
timestamp 1669390400
transform 1 0 5152 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_37
timestamp 1669390400
transform 1 0 5488 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_80_101
timestamp 1669390400
transform 1 0 12656 0 1 65856
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_105
timestamp 1669390400
transform 1 0 13104 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_108
timestamp 1669390400
transform 1 0 13440 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_80_172
timestamp 1669390400
transform 1 0 20608 0 1 65856
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_176
timestamp 1669390400
transform 1 0 21056 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_179
timestamp 1669390400
transform 1 0 21392 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_80_243
timestamp 1669390400
transform 1 0 28560 0 1 65856
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_247
timestamp 1669390400
transform 1 0 29008 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_250
timestamp 1669390400
transform 1 0 29344 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_80_314
timestamp 1669390400
transform 1 0 36512 0 1 65856
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_318
timestamp 1669390400
transform 1 0 36960 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_321
timestamp 1669390400
transform 1 0 37296 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_80_385
timestamp 1669390400
transform 1 0 44464 0 1 65856
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_389
timestamp 1669390400
transform 1 0 44912 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_392
timestamp 1669390400
transform 1 0 45248 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_80_456
timestamp 1669390400
transform 1 0 52416 0 1 65856
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_460
timestamp 1669390400
transform 1 0 52864 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_463
timestamp 1669390400
transform 1 0 53200 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_80_527
timestamp 1669390400
transform 1 0 60368 0 1 65856
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_531
timestamp 1669390400
transform 1 0 60816 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_534
timestamp 1669390400
transform 1 0 61152 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_80_598
timestamp 1669390400
transform 1 0 68320 0 1 65856
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_602
timestamp 1669390400
transform 1 0 68768 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_605
timestamp 1669390400
transform 1 0 69104 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_80_669
timestamp 1669390400
transform 1 0 76272 0 1 65856
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_673
timestamp 1669390400
transform 1 0 76720 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_80_676
timestamp 1669390400
transform 1 0 77056 0 1 65856
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_80_684
timestamp 1669390400
transform 1 0 77952 0 1 65856
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_2
timestamp 1669390400
transform 1 0 1568 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_81_66
timestamp 1669390400
transform 1 0 8736 0 -1 67424
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_70
timestamp 1669390400
transform 1 0 9184 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_73
timestamp 1669390400
transform 1 0 9520 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_81_137
timestamp 1669390400
transform 1 0 16688 0 -1 67424
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_141
timestamp 1669390400
transform 1 0 17136 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_144
timestamp 1669390400
transform 1 0 17472 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_81_208
timestamp 1669390400
transform 1 0 24640 0 -1 67424
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_212
timestamp 1669390400
transform 1 0 25088 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_215
timestamp 1669390400
transform 1 0 25424 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_81_279
timestamp 1669390400
transform 1 0 32592 0 -1 67424
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_283
timestamp 1669390400
transform 1 0 33040 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_286
timestamp 1669390400
transform 1 0 33376 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_81_350
timestamp 1669390400
transform 1 0 40544 0 -1 67424
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_354
timestamp 1669390400
transform 1 0 40992 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_357
timestamp 1669390400
transform 1 0 41328 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_81_421
timestamp 1669390400
transform 1 0 48496 0 -1 67424
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_425
timestamp 1669390400
transform 1 0 48944 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_428
timestamp 1669390400
transform 1 0 49280 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_81_492
timestamp 1669390400
transform 1 0 56448 0 -1 67424
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_496
timestamp 1669390400
transform 1 0 56896 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_499
timestamp 1669390400
transform 1 0 57232 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_81_563
timestamp 1669390400
transform 1 0 64400 0 -1 67424
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_567
timestamp 1669390400
transform 1 0 64848 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_570
timestamp 1669390400
transform 1 0 65184 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_81_634
timestamp 1669390400
transform 1 0 72352 0 -1 67424
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_638
timestamp 1669390400
transform 1 0 72800 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_81_641
timestamp 1669390400
transform 1 0 73136 0 -1 67424
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_81_673
timestamp 1669390400
transform 1 0 76720 0 -1 67424
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_81_681
timestamp 1669390400
transform 1 0 77616 0 -1 67424
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_685
timestamp 1669390400
transform 1 0 78064 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_687
timestamp 1669390400
transform 1 0 78288 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_82_2
timestamp 1669390400
transform 1 0 1568 0 1 67424
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_34
timestamp 1669390400
transform 1 0 5152 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_37
timestamp 1669390400
transform 1 0 5488 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_82_101
timestamp 1669390400
transform 1 0 12656 0 1 67424
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_105
timestamp 1669390400
transform 1 0 13104 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_108
timestamp 1669390400
transform 1 0 13440 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_82_172
timestamp 1669390400
transform 1 0 20608 0 1 67424
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_176
timestamp 1669390400
transform 1 0 21056 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_179
timestamp 1669390400
transform 1 0 21392 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_82_243
timestamp 1669390400
transform 1 0 28560 0 1 67424
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_247
timestamp 1669390400
transform 1 0 29008 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_250
timestamp 1669390400
transform 1 0 29344 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_82_314
timestamp 1669390400
transform 1 0 36512 0 1 67424
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_318
timestamp 1669390400
transform 1 0 36960 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_321
timestamp 1669390400
transform 1 0 37296 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_82_385
timestamp 1669390400
transform 1 0 44464 0 1 67424
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_389
timestamp 1669390400
transform 1 0 44912 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_392
timestamp 1669390400
transform 1 0 45248 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_82_456
timestamp 1669390400
transform 1 0 52416 0 1 67424
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_460
timestamp 1669390400
transform 1 0 52864 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_463
timestamp 1669390400
transform 1 0 53200 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_82_527
timestamp 1669390400
transform 1 0 60368 0 1 67424
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_531
timestamp 1669390400
transform 1 0 60816 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_534
timestamp 1669390400
transform 1 0 61152 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_82_598
timestamp 1669390400
transform 1 0 68320 0 1 67424
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_602
timestamp 1669390400
transform 1 0 68768 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_605
timestamp 1669390400
transform 1 0 69104 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_82_669
timestamp 1669390400
transform 1 0 76272 0 1 67424
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_673
timestamp 1669390400
transform 1 0 76720 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_82_676
timestamp 1669390400
transform 1 0 77056 0 1 67424
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_82_684
timestamp 1669390400
transform 1 0 77952 0 1 67424
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_2
timestamp 1669390400
transform 1 0 1568 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_83_66
timestamp 1669390400
transform 1 0 8736 0 -1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_70
timestamp 1669390400
transform 1 0 9184 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_73
timestamp 1669390400
transform 1 0 9520 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_83_137
timestamp 1669390400
transform 1 0 16688 0 -1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_141
timestamp 1669390400
transform 1 0 17136 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_144
timestamp 1669390400
transform 1 0 17472 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_83_208
timestamp 1669390400
transform 1 0 24640 0 -1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_212
timestamp 1669390400
transform 1 0 25088 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_215
timestamp 1669390400
transform 1 0 25424 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_83_279
timestamp 1669390400
transform 1 0 32592 0 -1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_283
timestamp 1669390400
transform 1 0 33040 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_286
timestamp 1669390400
transform 1 0 33376 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_83_350
timestamp 1669390400
transform 1 0 40544 0 -1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_354
timestamp 1669390400
transform 1 0 40992 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_357
timestamp 1669390400
transform 1 0 41328 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_83_421
timestamp 1669390400
transform 1 0 48496 0 -1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_425
timestamp 1669390400
transform 1 0 48944 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_428
timestamp 1669390400
transform 1 0 49280 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_83_492
timestamp 1669390400
transform 1 0 56448 0 -1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_496
timestamp 1669390400
transform 1 0 56896 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_499
timestamp 1669390400
transform 1 0 57232 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_83_563
timestamp 1669390400
transform 1 0 64400 0 -1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_567
timestamp 1669390400
transform 1 0 64848 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_570
timestamp 1669390400
transform 1 0 65184 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_83_634
timestamp 1669390400
transform 1 0 72352 0 -1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_638
timestamp 1669390400
transform 1 0 72800 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_83_641
timestamp 1669390400
transform 1 0 73136 0 -1 68992
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_83_673
timestamp 1669390400
transform 1 0 76720 0 -1 68992
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_83_681
timestamp 1669390400
transform 1 0 77616 0 -1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_685
timestamp 1669390400
transform 1 0 78064 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_687
timestamp 1669390400
transform 1 0 78288 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_84_2
timestamp 1669390400
transform 1 0 1568 0 1 68992
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_34
timestamp 1669390400
transform 1 0 5152 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_37
timestamp 1669390400
transform 1 0 5488 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_84_101
timestamp 1669390400
transform 1 0 12656 0 1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_105
timestamp 1669390400
transform 1 0 13104 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_108
timestamp 1669390400
transform 1 0 13440 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_84_172
timestamp 1669390400
transform 1 0 20608 0 1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_176
timestamp 1669390400
transform 1 0 21056 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_179
timestamp 1669390400
transform 1 0 21392 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_84_243
timestamp 1669390400
transform 1 0 28560 0 1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_247
timestamp 1669390400
transform 1 0 29008 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_250
timestamp 1669390400
transform 1 0 29344 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_84_314
timestamp 1669390400
transform 1 0 36512 0 1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_318
timestamp 1669390400
transform 1 0 36960 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_16  FILLER_84_321
timestamp 1669390400
transform 1 0 37296 0 1 68992
box 0 -60 1792 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_84_337
timestamp 1669390400
transform 1 0 39088 0 1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_341
timestamp 1669390400
transform 1 0 39536 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_344
timestamp 1669390400
transform 1 0 39872 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_346
timestamp 1669390400
transform 1 0 40096 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_349
timestamp 1669390400
transform 1 0 40432 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_84_353
timestamp 1669390400
transform 1 0 40880 0 1 68992
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_84_385
timestamp 1669390400
transform 1 0 44464 0 1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_389
timestamp 1669390400
transform 1 0 44912 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_84_392
timestamp 1669390400
transform 1 0 45248 0 1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_396
timestamp 1669390400
transform 1 0 45696 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_398
timestamp 1669390400
transform 1 0 45920 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_401
timestamp 1669390400
transform 1 0 46256 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_84_405
timestamp 1669390400
transform 1 0 46704 0 1 68992
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_16  FILLER_84_437
timestamp 1669390400
transform 1 0 50288 0 1 68992
box 0 -60 1792 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_453
timestamp 1669390400
transform 1 0 52080 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_456
timestamp 1669390400
transform 1 0 52416 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_460
timestamp 1669390400
transform 1 0 52864 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_463
timestamp 1669390400
transform 1 0 53200 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_84_527
timestamp 1669390400
transform 1 0 60368 0 1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_531
timestamp 1669390400
transform 1 0 60816 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_534
timestamp 1669390400
transform 1 0 61152 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_84_598
timestamp 1669390400
transform 1 0 68320 0 1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_602
timestamp 1669390400
transform 1 0 68768 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_605
timestamp 1669390400
transform 1 0 69104 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_84_669
timestamp 1669390400
transform 1 0 76272 0 1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_673
timestamp 1669390400
transform 1 0 76720 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_84_676
timestamp 1669390400
transform 1 0 77056 0 1 68992
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_84_684
timestamp 1669390400
transform 1 0 77952 0 1 68992
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_2
timestamp 1669390400
transform 1 0 1568 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_85_66
timestamp 1669390400
transform 1 0 8736 0 -1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_70
timestamp 1669390400
transform 1 0 9184 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_73
timestamp 1669390400
transform 1 0 9520 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_85_137
timestamp 1669390400
transform 1 0 16688 0 -1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_141
timestamp 1669390400
transform 1 0 17136 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_144
timestamp 1669390400
transform 1 0 17472 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_85_208
timestamp 1669390400
transform 1 0 24640 0 -1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_212
timestamp 1669390400
transform 1 0 25088 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_215
timestamp 1669390400
transform 1 0 25424 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_85_279
timestamp 1669390400
transform 1 0 32592 0 -1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_283
timestamp 1669390400
transform 1 0 33040 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_85_286
timestamp 1669390400
transform 1 0 33376 0 -1 70560
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_320
timestamp 1669390400
transform 1 0 37184 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_324
timestamp 1669390400
transform 1 0 37632 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_328
timestamp 1669390400
transform 1 0 38080 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_332
timestamp 1669390400
transform 1 0 38528 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_338
timestamp 1669390400
transform 1 0 39200 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_344
timestamp 1669390400
transform 1 0 39872 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_350
timestamp 1669390400
transform 1 0 40544 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_354
timestamp 1669390400
transform 1 0 40992 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_357
timestamp 1669390400
transform 1 0 41328 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_85_362
timestamp 1669390400
transform 1 0 41888 0 -1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_374
timestamp 1669390400
transform 1 0 43232 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_384
timestamp 1669390400
transform 1 0 44352 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_388
timestamp 1669390400
transform 1 0 44800 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_392
timestamp 1669390400
transform 1 0 45248 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_85_396
timestamp 1669390400
transform 1 0 45696 0 -1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_400
timestamp 1669390400
transform 1 0 46144 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_403
timestamp 1669390400
transform 1 0 46480 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_407
timestamp 1669390400
transform 1 0 46928 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_85_411
timestamp 1669390400
transform 1 0 47376 0 -1 70560
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_85_421
timestamp 1669390400
transform 1 0 48496 0 -1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_425
timestamp 1669390400
transform 1 0 48944 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_85_428
timestamp 1669390400
transform 1 0 49280 0 -1 70560
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_436
timestamp 1669390400
transform 1 0 50176 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_85_439
timestamp 1669390400
transform 1 0 50512 0 -1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_443
timestamp 1669390400
transform 1 0 50960 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_447
timestamp 1669390400
transform 1 0 51408 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_451
timestamp 1669390400
transform 1 0 51856 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_455
timestamp 1669390400
transform 1 0 52304 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_459
timestamp 1669390400
transform 1 0 52752 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_463
timestamp 1669390400
transform 1 0 53200 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_85_467
timestamp 1669390400
transform 1 0 53648 0 -1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_471
timestamp 1669390400
transform 1 0 54096 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_473
timestamp 1669390400
transform 1 0 54320 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_476
timestamp 1669390400
transform 1 0 54656 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_480
timestamp 1669390400
transform 1 0 55104 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_85_484
timestamp 1669390400
transform 1 0 55552 0 -1 70560
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_85_492
timestamp 1669390400
transform 1 0 56448 0 -1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_496
timestamp 1669390400
transform 1 0 56896 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_499
timestamp 1669390400
transform 1 0 57232 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_85_563
timestamp 1669390400
transform 1 0 64400 0 -1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_567
timestamp 1669390400
transform 1 0 64848 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_570
timestamp 1669390400
transform 1 0 65184 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_85_634
timestamp 1669390400
transform 1 0 72352 0 -1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_638
timestamp 1669390400
transform 1 0 72800 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_85_641
timestamp 1669390400
transform 1 0 73136 0 -1 70560
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_85_673
timestamp 1669390400
transform 1 0 76720 0 -1 70560
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_85_681
timestamp 1669390400
transform 1 0 77616 0 -1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_685
timestamp 1669390400
transform 1 0 78064 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_687
timestamp 1669390400
transform 1 0 78288 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_86_2
timestamp 1669390400
transform 1 0 1568 0 1 70560
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_34
timestamp 1669390400
transform 1 0 5152 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_37
timestamp 1669390400
transform 1 0 5488 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_86_101
timestamp 1669390400
transform 1 0 12656 0 1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_105
timestamp 1669390400
transform 1 0 13104 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_108
timestamp 1669390400
transform 1 0 13440 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_86_172
timestamp 1669390400
transform 1 0 20608 0 1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_176
timestamp 1669390400
transform 1 0 21056 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_179
timestamp 1669390400
transform 1 0 21392 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_86_243
timestamp 1669390400
transform 1 0 28560 0 1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_247
timestamp 1669390400
transform 1 0 29008 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_86_250
timestamp 1669390400
transform 1 0 29344 0 1 70560
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_86_282
timestamp 1669390400
transform 1 0 32928 0 1 70560
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_86_290
timestamp 1669390400
transform 1 0 33824 0 1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_294
timestamp 1669390400
transform 1 0 34272 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_296
timestamp 1669390400
transform 1 0 34496 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_299
timestamp 1669390400
transform 1 0 34832 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_301
timestamp 1669390400
transform 1 0 35056 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_86_304
timestamp 1669390400
transform 1 0 35392 0 1 70560
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_314
timestamp 1669390400
transform 1 0 36512 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_318
timestamp 1669390400
transform 1 0 36960 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_321
timestamp 1669390400
transform 1 0 37296 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_325
timestamp 1669390400
transform 1 0 37744 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_329
timestamp 1669390400
transform 1 0 38192 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_339
timestamp 1669390400
transform 1 0 39312 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_347
timestamp 1669390400
transform 1 0 40208 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_349
timestamp 1669390400
transform 1 0 40432 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_363
timestamp 1669390400
transform 1 0 42000 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_389
timestamp 1669390400
transform 1 0 44912 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_392
timestamp 1669390400
transform 1 0 45248 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_395
timestamp 1669390400
transform 1 0 45584 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_399
timestamp 1669390400
transform 1 0 46032 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_403
timestamp 1669390400
transform 1 0 46480 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_86_407
timestamp 1669390400
transform 1 0 46928 0 1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_413
timestamp 1669390400
transform 1 0 47600 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_417
timestamp 1669390400
transform 1 0 48048 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_421
timestamp 1669390400
transform 1 0 48496 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_425
timestamp 1669390400
transform 1 0 48944 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_429
timestamp 1669390400
transform 1 0 49392 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_86_433
timestamp 1669390400
transform 1 0 49840 0 1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_439
timestamp 1669390400
transform 1 0 50512 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_86_443
timestamp 1669390400
transform 1 0 50960 0 1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_451
timestamp 1669390400
transform 1 0 51856 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_86_457
timestamp 1669390400
transform 1 0 52528 0 1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_463
timestamp 1669390400
transform 1 0 53200 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_469
timestamp 1669390400
transform 1 0 53872 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_473
timestamp 1669390400
transform 1 0 54320 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_475
timestamp 1669390400
transform 1 0 54544 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_478
timestamp 1669390400
transform 1 0 54880 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_480
timestamp 1669390400
transform 1 0 55104 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_483
timestamp 1669390400
transform 1 0 55440 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_487
timestamp 1669390400
transform 1 0 55888 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_512
timestamp 1669390400
transform 1 0 58688 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_16  FILLER_86_516
timestamp 1669390400
transform 1 0 59136 0 1 70560
box 0 -60 1792 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_534
timestamp 1669390400
transform 1 0 61152 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_86_598
timestamp 1669390400
transform 1 0 68320 0 1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_602
timestamp 1669390400
transform 1 0 68768 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_605
timestamp 1669390400
transform 1 0 69104 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_86_669
timestamp 1669390400
transform 1 0 76272 0 1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_673
timestamp 1669390400
transform 1 0 76720 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_86_676
timestamp 1669390400
transform 1 0 77056 0 1 70560
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_86_684
timestamp 1669390400
transform 1 0 77952 0 1 70560
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_2
timestamp 1669390400
transform 1 0 1568 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_87_66
timestamp 1669390400
transform 1 0 8736 0 -1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_70
timestamp 1669390400
transform 1 0 9184 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_73
timestamp 1669390400
transform 1 0 9520 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_87_137
timestamp 1669390400
transform 1 0 16688 0 -1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_141
timestamp 1669390400
transform 1 0 17136 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_144
timestamp 1669390400
transform 1 0 17472 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_87_208
timestamp 1669390400
transform 1 0 24640 0 -1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_212
timestamp 1669390400
transform 1 0 25088 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_215
timestamp 1669390400
transform 1 0 25424 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_87_279
timestamp 1669390400
transform 1 0 32592 0 -1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_283
timestamp 1669390400
transform 1 0 33040 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_87_286
timestamp 1669390400
transform 1 0 33376 0 -1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_292
timestamp 1669390400
transform 1 0 34048 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_296
timestamp 1669390400
transform 1 0 34496 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_300
timestamp 1669390400
transform 1 0 34944 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_302
timestamp 1669390400
transform 1 0 35168 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_307
timestamp 1669390400
transform 1 0 35728 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_311
timestamp 1669390400
transform 1 0 36176 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_315
timestamp 1669390400
transform 1 0 36624 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_321
timestamp 1669390400
transform 1 0 37296 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_329
timestamp 1669390400
transform 1 0 38192 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_354
timestamp 1669390400
transform 1 0 40992 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_357
timestamp 1669390400
transform 1 0 41328 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_360
timestamp 1669390400
transform 1 0 41664 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_87_385
timestamp 1669390400
transform 1 0 44464 0 -1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_394
timestamp 1669390400
transform 1 0 45472 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_401
timestamp 1669390400
transform 1 0 46256 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_407
timestamp 1669390400
transform 1 0 46928 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_411
timestamp 1669390400
transform 1 0 47376 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_415
timestamp 1669390400
transform 1 0 47824 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_419
timestamp 1669390400
transform 1 0 48272 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_423
timestamp 1669390400
transform 1 0 48720 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_425
timestamp 1669390400
transform 1 0 48944 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_428
timestamp 1669390400
transform 1 0 49280 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_453
timestamp 1669390400
transform 1 0 52080 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_87_463
timestamp 1669390400
transform 1 0 53200 0 -1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_467
timestamp 1669390400
transform 1 0 53648 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_476
timestamp 1669390400
transform 1 0 54656 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_478
timestamp 1669390400
transform 1 0 54880 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_485
timestamp 1669390400
transform 1 0 55664 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_495
timestamp 1669390400
transform 1 0 56784 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_499
timestamp 1669390400
transform 1 0 57232 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_513
timestamp 1669390400
transform 1 0 58800 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_517
timestamp 1669390400
transform 1 0 59248 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_87_521
timestamp 1669390400
transform 1 0 59696 0 -1 72128
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_87_553
timestamp 1669390400
transform 1 0 63280 0 -1 72128
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_87_561
timestamp 1669390400
transform 1 0 64176 0 -1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_565
timestamp 1669390400
transform 1 0 64624 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_567
timestamp 1669390400
transform 1 0 64848 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_570
timestamp 1669390400
transform 1 0 65184 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_87_634
timestamp 1669390400
transform 1 0 72352 0 -1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_638
timestamp 1669390400
transform 1 0 72800 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_87_641
timestamp 1669390400
transform 1 0 73136 0 -1 72128
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_87_673
timestamp 1669390400
transform 1 0 76720 0 -1 72128
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_87_681
timestamp 1669390400
transform 1 0 77616 0 -1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_685
timestamp 1669390400
transform 1 0 78064 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_687
timestamp 1669390400
transform 1 0 78288 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_88_2
timestamp 1669390400
transform 1 0 1568 0 1 72128
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_34
timestamp 1669390400
transform 1 0 5152 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_37
timestamp 1669390400
transform 1 0 5488 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_88_101
timestamp 1669390400
transform 1 0 12656 0 1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_105
timestamp 1669390400
transform 1 0 13104 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_108
timestamp 1669390400
transform 1 0 13440 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_88_172
timestamp 1669390400
transform 1 0 20608 0 1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_176
timestamp 1669390400
transform 1 0 21056 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_179
timestamp 1669390400
transform 1 0 21392 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_88_243
timestamp 1669390400
transform 1 0 28560 0 1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_247
timestamp 1669390400
transform 1 0 29008 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_88_250
timestamp 1669390400
transform 1 0 29344 0 1 72128
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_88_258
timestamp 1669390400
transform 1 0 30240 0 1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_262
timestamp 1669390400
transform 1 0 30688 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_88_265
timestamp 1669390400
transform 1 0 31024 0 1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_269
timestamp 1669390400
transform 1 0 31472 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_271
timestamp 1669390400
transform 1 0 31696 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_88_274
timestamp 1669390400
transform 1 0 32032 0 1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_280
timestamp 1669390400
transform 1 0 32704 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_284
timestamp 1669390400
transform 1 0 33152 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_288
timestamp 1669390400
transform 1 0 33600 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_292
timestamp 1669390400
transform 1 0 34048 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_298
timestamp 1669390400
transform 1 0 34720 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_304
timestamp 1669390400
transform 1 0 35392 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_306
timestamp 1669390400
transform 1 0 35616 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_311
timestamp 1669390400
transform 1 0 36176 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_318
timestamp 1669390400
transform 1 0 36960 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_321
timestamp 1669390400
transform 1 0 37296 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_327
timestamp 1669390400
transform 1 0 37968 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_88_352
timestamp 1669390400
transform 1 0 40768 0 1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_362
timestamp 1669390400
transform 1 0 41888 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_376
timestamp 1669390400
transform 1 0 43456 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_88_386
timestamp 1669390400
transform 1 0 44576 0 1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_392
timestamp 1669390400
transform 1 0 45248 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_405
timestamp 1669390400
transform 1 0 46704 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_411
timestamp 1669390400
transform 1 0 47376 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_417
timestamp 1669390400
transform 1 0 48048 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_423
timestamp 1669390400
transform 1 0 48720 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_425
timestamp 1669390400
transform 1 0 48944 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_430
timestamp 1669390400
transform 1 0 49504 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_440
timestamp 1669390400
transform 1 0 50624 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_444
timestamp 1669390400
transform 1 0 51072 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_446
timestamp 1669390400
transform 1 0 51296 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_460
timestamp 1669390400
transform 1 0 52864 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_463
timestamp 1669390400
transform 1 0 53200 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_476
timestamp 1669390400
transform 1 0 54656 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_484
timestamp 1669390400
transform 1 0 55552 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_488
timestamp 1669390400
transform 1 0 56000 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_490
timestamp 1669390400
transform 1 0 56224 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_514
timestamp 1669390400
transform 1 0 58912 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_520
timestamp 1669390400
transform 1 0 59584 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_524
timestamp 1669390400
transform 1 0 60032 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_88_528
timestamp 1669390400
transform 1 0 60480 0 1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_534
timestamp 1669390400
transform 1 0 61152 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_537
timestamp 1669390400
transform 1 0 61488 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_601
timestamp 1669390400
transform 1 0 68656 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_605
timestamp 1669390400
transform 1 0 69104 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_88_669
timestamp 1669390400
transform 1 0 76272 0 1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_673
timestamp 1669390400
transform 1 0 76720 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_88_676
timestamp 1669390400
transform 1 0 77056 0 1 72128
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_88_684
timestamp 1669390400
transform 1 0 77952 0 1 72128
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_2
timestamp 1669390400
transform 1 0 1568 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_89_66
timestamp 1669390400
transform 1 0 8736 0 -1 73696
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_70
timestamp 1669390400
transform 1 0 9184 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_73
timestamp 1669390400
transform 1 0 9520 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_89_137
timestamp 1669390400
transform 1 0 16688 0 -1 73696
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_141
timestamp 1669390400
transform 1 0 17136 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_144
timestamp 1669390400
transform 1 0 17472 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_89_208
timestamp 1669390400
transform 1 0 24640 0 -1 73696
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_212
timestamp 1669390400
transform 1 0 25088 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_89_215
timestamp 1669390400
transform 1 0 25424 0 -1 73696
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_247
timestamp 1669390400
transform 1 0 29008 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_249
timestamp 1669390400
transform 1 0 29232 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_252
timestamp 1669390400
transform 1 0 29568 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_256
timestamp 1669390400
transform 1 0 30016 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_262
timestamp 1669390400
transform 1 0 30688 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_264
timestamp 1669390400
transform 1 0 30912 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_271
timestamp 1669390400
transform 1 0 31696 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_89_277
timestamp 1669390400
transform 1 0 32368 0 -1 73696
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_283
timestamp 1669390400
transform 1 0 33040 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_286
timestamp 1669390400
transform 1 0 33376 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_293
timestamp 1669390400
transform 1 0 34160 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_89_301
timestamp 1669390400
transform 1 0 35056 0 -1 73696
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_309
timestamp 1669390400
transform 1 0 35952 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_326
timestamp 1669390400
transform 1 0 37856 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_340
timestamp 1669390400
transform 1 0 39424 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_342
timestamp 1669390400
transform 1 0 39648 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_345
timestamp 1669390400
transform 1 0 39984 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_354
timestamp 1669390400
transform 1 0 40992 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_357
timestamp 1669390400
transform 1 0 41328 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_89_363
timestamp 1669390400
transform 1 0 42000 0 -1 73696
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_377
timestamp 1669390400
transform 1 0 43568 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_381
timestamp 1669390400
transform 1 0 44016 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_383
timestamp 1669390400
transform 1 0 44240 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_395
timestamp 1669390400
transform 1 0 45584 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_409
timestamp 1669390400
transform 1 0 47152 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_89_415
timestamp 1669390400
transform 1 0 47824 0 -1 73696
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_425
timestamp 1669390400
transform 1 0 48944 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_428
timestamp 1669390400
transform 1 0 49280 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_440
timestamp 1669390400
transform 1 0 50624 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_446
timestamp 1669390400
transform 1 0 51296 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_471
timestamp 1669390400
transform 1 0 54096 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_481
timestamp 1669390400
transform 1 0 55216 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_485
timestamp 1669390400
transform 1 0 55664 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_495
timestamp 1669390400
transform 1 0 56784 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_499
timestamp 1669390400
transform 1 0 57232 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_89_506
timestamp 1669390400
transform 1 0 58016 0 -1 73696
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_522
timestamp 1669390400
transform 1 0 59808 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_528
timestamp 1669390400
transform 1 0 60480 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_534
timestamp 1669390400
transform 1 0 61152 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_538
timestamp 1669390400
transform 1 0 61600 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_542
timestamp 1669390400
transform 1 0 62048 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_546
timestamp 1669390400
transform 1 0 62496 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_16  FILLER_89_550
timestamp 1669390400
transform 1 0 62944 0 -1 73696
box 0 -60 1792 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_566
timestamp 1669390400
transform 1 0 64736 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_570
timestamp 1669390400
transform 1 0 65184 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_89_634
timestamp 1669390400
transform 1 0 72352 0 -1 73696
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_638
timestamp 1669390400
transform 1 0 72800 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_89_641
timestamp 1669390400
transform 1 0 73136 0 -1 73696
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_89_673
timestamp 1669390400
transform 1 0 76720 0 -1 73696
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_89_681
timestamp 1669390400
transform 1 0 77616 0 -1 73696
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_685
timestamp 1669390400
transform 1 0 78064 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_687
timestamp 1669390400
transform 1 0 78288 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_90_2
timestamp 1669390400
transform 1 0 1568 0 1 73696
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_34
timestamp 1669390400
transform 1 0 5152 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_37
timestamp 1669390400
transform 1 0 5488 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_90_101
timestamp 1669390400
transform 1 0 12656 0 1 73696
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_105
timestamp 1669390400
transform 1 0 13104 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_108
timestamp 1669390400
transform 1 0 13440 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_90_172
timestamp 1669390400
transform 1 0 20608 0 1 73696
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_176
timestamp 1669390400
transform 1 0 21056 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_179
timestamp 1669390400
transform 1 0 21392 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_243
timestamp 1669390400
transform 1 0 28560 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_247
timestamp 1669390400
transform 1 0 29008 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_250
timestamp 1669390400
transform 1 0 29344 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_254
timestamp 1669390400
transform 1 0 29792 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_262
timestamp 1669390400
transform 1 0 30688 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_270
timestamp 1669390400
transform 1 0 31584 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_278
timestamp 1669390400
transform 1 0 32480 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_90_288
timestamp 1669390400
transform 1 0 33600 0 1 73696
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_300
timestamp 1669390400
transform 1 0 34944 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_310
timestamp 1669390400
transform 1 0 36064 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_312
timestamp 1669390400
transform 1 0 36288 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_318
timestamp 1669390400
transform 1 0 36960 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_321
timestamp 1669390400
transform 1 0 37296 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_332
timestamp 1669390400
transform 1 0 38528 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_342
timestamp 1669390400
transform 1 0 39648 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_344
timestamp 1669390400
transform 1 0 39872 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_347
timestamp 1669390400
transform 1 0 40208 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_357
timestamp 1669390400
transform 1 0 41328 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_359
timestamp 1669390400
transform 1 0 41552 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_377
timestamp 1669390400
transform 1 0 43568 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_387
timestamp 1669390400
transform 1 0 44688 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_389
timestamp 1669390400
transform 1 0 44912 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_392
timestamp 1669390400
transform 1 0 45248 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_394
timestamp 1669390400
transform 1 0 45472 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_405
timestamp 1669390400
transform 1 0 46704 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_411
timestamp 1669390400
transform 1 0 47376 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_417
timestamp 1669390400
transform 1 0 48048 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_423
timestamp 1669390400
transform 1 0 48720 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_429
timestamp 1669390400
transform 1 0 49392 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_441
timestamp 1669390400
transform 1 0 50736 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_452
timestamp 1669390400
transform 1 0 51968 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_459
timestamp 1669390400
transform 1 0 52752 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_463
timestamp 1669390400
transform 1 0 53200 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_481
timestamp 1669390400
transform 1 0 55216 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_493
timestamp 1669390400
transform 1 0 56560 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_495
timestamp 1669390400
transform 1 0 56784 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_502
timestamp 1669390400
transform 1 0 57568 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_90_509
timestamp 1669390400
transform 1 0 58352 0 1 73696
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_513
timestamp 1669390400
transform 1 0 58800 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_524
timestamp 1669390400
transform 1 0 60032 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_531
timestamp 1669390400
transform 1 0 60816 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_534
timestamp 1669390400
transform 1 0 61152 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_539
timestamp 1669390400
transform 1 0 61712 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_543
timestamp 1669390400
transform 1 0 62160 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_547
timestamp 1669390400
transform 1 0 62608 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_551
timestamp 1669390400
transform 1 0 63056 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_90_555
timestamp 1669390400
transform 1 0 63504 0 1 73696
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_16  FILLER_90_587
timestamp 1669390400
transform 1 0 67088 0 1 73696
box 0 -60 1792 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_605
timestamp 1669390400
transform 1 0 69104 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_90_669
timestamp 1669390400
transform 1 0 76272 0 1 73696
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_673
timestamp 1669390400
transform 1 0 76720 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_90_676
timestamp 1669390400
transform 1 0 77056 0 1 73696
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_684
timestamp 1669390400
transform 1 0 77952 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_687
timestamp 1669390400
transform 1 0 78288 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_2
timestamp 1669390400
transform 1 0 1568 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_91_66
timestamp 1669390400
transform 1 0 8736 0 -1 75264
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_70
timestamp 1669390400
transform 1 0 9184 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_73
timestamp 1669390400
transform 1 0 9520 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_91_137
timestamp 1669390400
transform 1 0 16688 0 -1 75264
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_141
timestamp 1669390400
transform 1 0 17136 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_144
timestamp 1669390400
transform 1 0 17472 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_91_208
timestamp 1669390400
transform 1 0 24640 0 -1 75264
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_212
timestamp 1669390400
transform 1 0 25088 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_16  FILLER_91_215
timestamp 1669390400
transform 1 0 25424 0 -1 75264
box 0 -60 1792 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_91_231
timestamp 1669390400
transform 1 0 27216 0 -1 75264
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_235
timestamp 1669390400
transform 1 0 27664 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_237
timestamp 1669390400
transform 1 0 27888 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_240
timestamp 1669390400
transform 1 0 28224 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_244
timestamp 1669390400
transform 1 0 28672 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_252
timestamp 1669390400
transform 1 0 29568 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_260
timestamp 1669390400
transform 1 0 30464 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_91_270
timestamp 1669390400
transform 1 0 31584 0 -1 75264
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_274
timestamp 1669390400
transform 1 0 32032 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_283
timestamp 1669390400
transform 1 0 33040 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_286
timestamp 1669390400
transform 1 0 33376 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_290
timestamp 1669390400
transform 1 0 33824 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_300
timestamp 1669390400
transform 1 0 34944 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_310
timestamp 1669390400
transform 1 0 36064 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_327
timestamp 1669390400
transform 1 0 37968 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_329
timestamp 1669390400
transform 1 0 38192 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_336
timestamp 1669390400
transform 1 0 38976 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_346
timestamp 1669390400
transform 1 0 40096 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_354
timestamp 1669390400
transform 1 0 40992 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_357
timestamp 1669390400
transform 1 0 41328 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_91_364
timestamp 1669390400
transform 1 0 42112 0 -1 75264
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_378
timestamp 1669390400
transform 1 0 43680 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_91_389
timestamp 1669390400
transform 1 0 44912 0 -1 75264
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_401
timestamp 1669390400
transform 1 0 46256 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_408
timestamp 1669390400
transform 1 0 47040 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_425
timestamp 1669390400
transform 1 0 48944 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_428
timestamp 1669390400
transform 1 0 49280 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_91_439
timestamp 1669390400
transform 1 0 50512 0 -1 75264
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_443
timestamp 1669390400
transform 1 0 50960 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_91_456
timestamp 1669390400
transform 1 0 52416 0 -1 75264
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_466
timestamp 1669390400
transform 1 0 53536 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_478
timestamp 1669390400
transform 1 0 54880 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_488
timestamp 1669390400
transform 1 0 56000 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_496
timestamp 1669390400
transform 1 0 56896 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_499
timestamp 1669390400
transform 1 0 57232 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_515
timestamp 1669390400
transform 1 0 59024 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_525
timestamp 1669390400
transform 1 0 60144 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_532
timestamp 1669390400
transform 1 0 60928 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_538
timestamp 1669390400
transform 1 0 61600 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_544
timestamp 1669390400
transform 1 0 62272 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_550
timestamp 1669390400
transform 1 0 62944 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_556
timestamp 1669390400
transform 1 0 63616 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_562
timestamp 1669390400
transform 1 0 64288 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_566
timestamp 1669390400
transform 1 0 64736 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_570
timestamp 1669390400
transform 1 0 65184 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_16  FILLER_91_573
timestamp 1669390400
transform 1 0 65520 0 -1 75264
box 0 -60 1792 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_91_589
timestamp 1669390400
transform 1 0 67312 0 -1 75264
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_601
timestamp 1669390400
transform 1 0 68656 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_603
timestamp 1669390400
transform 1 0 68880 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_91_606
timestamp 1669390400
transform 1 0 69216 0 -1 75264
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_91_614
timestamp 1669390400
transform 1 0 70112 0 -1 75264
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_618
timestamp 1669390400
transform 1 0 70560 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_16  FILLER_91_621
timestamp 1669390400
transform 1 0 70896 0 -1 75264
box 0 -60 1792 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_637
timestamp 1669390400
transform 1 0 72688 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_641
timestamp 1669390400
transform 1 0 73136 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_91_644
timestamp 1669390400
transform 1 0 73472 0 -1 75264
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_652
timestamp 1669390400
transform 1 0 74368 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_687
timestamp 1669390400
transform 1 0 78288 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_2
timestamp 1669390400
transform 1 0 1568 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_16  FILLER_92_5
timestamp 1669390400
transform 1 0 1904 0 1 75264
box 0 -60 1792 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_92_21
timestamp 1669390400
transform 1 0 3696 0 1 75264
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_92_29
timestamp 1669390400
transform 1 0 4592 0 1 75264
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_33
timestamp 1669390400
transform 1 0 5040 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_37
timestamp 1669390400
transform 1 0 5488 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_92_43
timestamp 1669390400
transform 1 0 6160 0 1 75264
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_55
timestamp 1669390400
transform 1 0 7504 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_32  FILLER_92_59
timestamp 1669390400
transform 1 0 7952 0 1 75264
box 0 -60 3584 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_92_91
timestamp 1669390400
transform 1 0 11536 0 1 75264
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_92_99
timestamp 1669390400
transform 1 0 12432 0 1 75264
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_105
timestamp 1669390400
transform 1 0 13104 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_108
timestamp 1669390400
transform 1 0 13440 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_92_113
timestamp 1669390400
transform 1 0 14000 0 1 75264
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_121
timestamp 1669390400
transform 1 0 14896 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_127
timestamp 1669390400
transform 1 0 15568 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_92_131
timestamp 1669390400
transform 1 0 16016 0 1 75264
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_139
timestamp 1669390400
transform 1 0 16912 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_145
timestamp 1669390400
transform 1 0 17584 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_92_149
timestamp 1669390400
transform 1 0 18032 0 1 75264
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_157
timestamp 1669390400
transform 1 0 18928 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_163
timestamp 1669390400
transform 1 0 19600 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_92_167
timestamp 1669390400
transform 1 0 20048 0 1 75264
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_171
timestamp 1669390400
transform 1 0 20496 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_173
timestamp 1669390400
transform 1 0 20720 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_176
timestamp 1669390400
transform 1 0 21056 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_179
timestamp 1669390400
transform 1 0 21392 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_92_184
timestamp 1669390400
transform 1 0 21952 0 1 75264
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_192
timestamp 1669390400
transform 1 0 22848 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_194
timestamp 1669390400
transform 1 0 23072 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_199
timestamp 1669390400
transform 1 0 23632 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_92_203
timestamp 1669390400
transform 1 0 24080 0 1 75264
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_207
timestamp 1669390400
transform 1 0 24528 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_211
timestamp 1669390400
transform 1 0 24976 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_8  FILLER_92_217
timestamp 1669390400
transform 1 0 25648 0 1 75264
box 0 -60 896 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_227
timestamp 1669390400
transform 1 0 26768 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_233
timestamp 1669390400
transform 1 0 27440 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_239
timestamp 1669390400
transform 1 0 28112 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_247
timestamp 1669390400
transform 1 0 29008 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_250
timestamp 1669390400
transform 1 0 29344 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_252
timestamp 1669390400
transform 1 0 29568 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_261
timestamp 1669390400
transform 1 0 30576 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_271
timestamp 1669390400
transform 1 0 31696 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_287
timestamp 1669390400
transform 1 0 33488 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_92_297
timestamp 1669390400
transform 1 0 34608 0 1 75264
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_307
timestamp 1669390400
transform 1 0 35728 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_318
timestamp 1669390400
transform 1 0 36960 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_321
timestamp 1669390400
transform 1 0 37296 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_325
timestamp 1669390400
transform 1 0 37744 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_341
timestamp 1669390400
transform 1 0 39536 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_353
timestamp 1669390400
transform 1 0 40880 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_355
timestamp 1669390400
transform 1 0 41104 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_358
timestamp 1669390400
transform 1 0 41440 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_366
timestamp 1669390400
transform 1 0 42336 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_378
timestamp 1669390400
transform 1 0 43680 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_92_386
timestamp 1669390400
transform 1 0 44576 0 1 75264
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_392
timestamp 1669390400
transform 1 0 45248 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_399
timestamp 1669390400
transform 1 0 46032 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_403
timestamp 1669390400
transform 1 0 46480 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_430
timestamp 1669390400
transform 1 0 49504 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_434
timestamp 1669390400
transform 1 0 49952 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_436
timestamp 1669390400
transform 1 0 50176 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_445
timestamp 1669390400
transform 1 0 51184 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_455
timestamp 1669390400
transform 1 0 52304 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_459
timestamp 1669390400
transform 1 0 52752 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_463
timestamp 1669390400
transform 1 0 53200 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_475
timestamp 1669390400
transform 1 0 54544 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_493
timestamp 1669390400
transform 1 0 56560 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_501
timestamp 1669390400
transform 1 0 57456 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_509
timestamp 1669390400
transform 1 0 58352 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_517
timestamp 1669390400
transform 1 0 59248 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_525
timestamp 1669390400
transform 1 0 60144 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_531
timestamp 1669390400
transform 1 0 60816 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_534
timestamp 1669390400
transform 1 0 61152 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_540
timestamp 1669390400
transform 1 0 61824 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_546
timestamp 1669390400
transform 1 0 62496 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_548
timestamp 1669390400
transform 1 0 62720 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_574
timestamp 1669390400
transform 1 0 65632 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_580
timestamp 1669390400
transform 1 0 66304 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_586
timestamp 1669390400
transform 1 0 66976 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_592
timestamp 1669390400
transform 1 0 67648 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_598
timestamp 1669390400
transform 1 0 68320 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_602
timestamp 1669390400
transform 1 0 68768 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_605
timestamp 1669390400
transform 1 0 69104 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_612
timestamp 1669390400
transform 1 0 69888 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_618
timestamp 1669390400
transform 1 0 70560 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_620
timestamp 1669390400
transform 1 0 70784 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_646
timestamp 1669390400
transform 1 0 73696 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_673
timestamp 1669390400
transform 1 0 76720 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_676
timestamp 1669390400
transform 1 0 77056 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_92_679
timestamp 1669390400
transform 1 0 77392 0 1 75264
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_687
timestamp 1669390400
transform 1 0 78288 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_2
timestamp 1669390400
transform 1 0 1568 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_19
timestamp 1669390400
transform 1 0 3472 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_93_25
timestamp 1669390400
transform 1 0 4144 0 -1 76832
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_29
timestamp 1669390400
transform 1 0 4592 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_34
timestamp 1669390400
transform 1 0 5152 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_37
timestamp 1669390400
transform 1 0 5488 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_93_52
timestamp 1669390400
transform 1 0 7168 0 -1 76832
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_56
timestamp 1669390400
transform 1 0 7616 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_93_61
timestamp 1669390400
transform 1 0 8176 0 -1 76832
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_69
timestamp 1669390400
transform 1 0 9072 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_72
timestamp 1669390400
transform 1 0 9408 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_74
timestamp 1669390400
transform 1 0 9632 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_93_79
timestamp 1669390400
transform 1 0 10192 0 -1 76832
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_83
timestamp 1669390400
transform 1 0 10640 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_88
timestamp 1669390400
transform 1 0 11200 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_104
timestamp 1669390400
transform 1 0 12992 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_107
timestamp 1669390400
transform 1 0 13328 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_123
timestamp 1669390400
transform 1 0 15120 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_139
timestamp 1669390400
transform 1 0 16912 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_142
timestamp 1669390400
transform 1 0 17248 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_158
timestamp 1669390400
transform 1 0 19040 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_174
timestamp 1669390400
transform 1 0 20832 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_177
timestamp 1669390400
transform 1 0 21168 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_193
timestamp 1669390400
transform 1 0 22960 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_209
timestamp 1669390400
transform 1 0 24752 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_212
timestamp 1669390400
transform 1 0 25088 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_228
timestamp 1669390400
transform 1 0 26880 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_244
timestamp 1669390400
transform 1 0 28672 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_247
timestamp 1669390400
transform 1 0 29008 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_253
timestamp 1669390400
transform 1 0 29680 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_93_269
timestamp 1669390400
transform 1 0 31472 0 -1 76832
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_279
timestamp 1669390400
transform 1 0 32592 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_282
timestamp 1669390400
transform 1 0 32928 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_298
timestamp 1669390400
transform 1 0 34720 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_314
timestamp 1669390400
transform 1 0 36512 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_317
timestamp 1669390400
transform 1 0 36848 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_323
timestamp 1669390400
transform 1 0 37520 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_331
timestamp 1669390400
transform 1 0 38416 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_349
timestamp 1669390400
transform 1 0 40432 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_352
timestamp 1669390400
transform 1 0 40768 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_369
timestamp 1669390400
transform 1 0 42672 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_380
timestamp 1669390400
transform 1 0 43904 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_384
timestamp 1669390400
transform 1 0 44352 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_387
timestamp 1669390400
transform 1 0 44688 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_394
timestamp 1669390400
transform 1 0 45472 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_402
timestamp 1669390400
transform 1 0 46368 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_410
timestamp 1669390400
transform 1 0 47264 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_412
timestamp 1669390400
transform 1 0 47488 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_419
timestamp 1669390400
transform 1 0 48272 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_422
timestamp 1669390400
transform 1 0 48608 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_428
timestamp 1669390400
transform 1 0 49280 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_93_437
timestamp 1669390400
transform 1 0 50288 0 -1 76832
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_446
timestamp 1669390400
transform 1 0 51296 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_454
timestamp 1669390400
transform 1 0 52192 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_457
timestamp 1669390400
transform 1 0 52528 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_483
timestamp 1669390400
transform 1 0 55440 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_489
timestamp 1669390400
transform 1 0 56112 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_492
timestamp 1669390400
transform 1 0 56448 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_494
timestamp 1669390400
transform 1 0 56672 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_511
timestamp 1669390400
transform 1 0 58576 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_519
timestamp 1669390400
transform 1 0 59472 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_523
timestamp 1669390400
transform 1 0 59920 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_4  FILLER_93_527
timestamp 1669390400
transform 1 0 60368 0 -1 76832
box 0 -60 448 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_537
timestamp 1669390400
transform 1 0 61488 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_543
timestamp 1669390400
transform 1 0 62160 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_549
timestamp 1669390400
transform 1 0 62832 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_555
timestamp 1669390400
transform 1 0 63504 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_559
timestamp 1669390400
transform 1 0 63952 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_562
timestamp 1669390400
transform 1 0 64288 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_565
timestamp 1669390400
transform 1 0 64624 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_592
timestamp 1669390400
transform 1 0 67648 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_594
timestamp 1669390400
transform 1 0 67872 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_597
timestamp 1669390400
transform 1 0 68208 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_623
timestamp 1669390400
transform 1 0 71120 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_629
timestamp 1669390400
transform 1 0 71792 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_632
timestamp 1669390400
transform 1 0 72128 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_637
timestamp 1669390400
transform 1 0 72688 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_645
timestamp 1669390400
transform 1 0 73584 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_651
timestamp 1669390400
transform 1 0 74256 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_657
timestamp 1669390400
transform 1 0 74928 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_663
timestamp 1669390400
transform 1 0 75600 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_667
timestamp 1669390400
transform 1 0 76048 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_672
timestamp 1669390400
transform 1 0 76608 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_678
timestamp 1669390400
transform 1 0 77280 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_680
timestamp 1669390400
transform 1 0 77504 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_685
timestamp 1669390400
transform 1 0 78064 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_687
timestamp 1669390400
transform 1 0 78288 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 78624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 78624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 78624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 78624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 78624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 78624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 78624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 78624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 78624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 78624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 78624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 78624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1669390400
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1669390400
transform -1 0 78624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1669390400
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1669390400
transform -1 0 78624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1669390400
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1669390400
transform -1 0 78624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1669390400
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1669390400
transform -1 0 78624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1669390400
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1669390400
transform -1 0 78624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1669390400
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1669390400
transform -1 0 78624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1669390400
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1669390400
transform -1 0 78624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1669390400
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1669390400
transform -1 0 78624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1669390400
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1669390400
transform -1 0 78624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1669390400
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1669390400
transform -1 0 78624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1669390400
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1669390400
transform -1 0 78624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1669390400
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1669390400
transform -1 0 78624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1669390400
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1669390400
transform -1 0 78624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1669390400
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1669390400
transform -1 0 78624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1669390400
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1669390400
transform -1 0 78624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1669390400
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1669390400
transform -1 0 78624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1669390400
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1669390400
transform -1 0 78624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1669390400
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1669390400
transform -1 0 78624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1669390400
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1669390400
transform -1 0 78624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1669390400
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1669390400
transform -1 0 78624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1669390400
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1669390400
transform -1 0 78624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1669390400
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1669390400
transform -1 0 78624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1669390400
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1669390400
transform -1 0 78624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1669390400
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1669390400
transform -1 0 78624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1669390400
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1669390400
transform -1 0 78624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1669390400
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1669390400
transform -1 0 78624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1669390400
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1669390400
transform -1 0 78624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1669390400
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1669390400
transform -1 0 78624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1669390400
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1669390400
transform -1 0 78624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1669390400
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1669390400
transform -1 0 78624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1669390400
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1669390400
transform -1 0 78624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1669390400
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1669390400
transform -1 0 78624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1669390400
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1669390400
transform -1 0 78624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1669390400
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1669390400
transform -1 0 78624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1669390400
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1669390400
transform -1 0 78624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1669390400
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1669390400
transform -1 0 78624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1669390400
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1669390400
transform -1 0 78624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1669390400
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1669390400
transform -1 0 78624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1669390400
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1669390400
transform -1 0 78624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1669390400
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1669390400
transform -1 0 78624 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1669390400
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1669390400
transform -1 0 78624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1669390400
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1669390400
transform -1 0 78624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1669390400
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1669390400
transform -1 0 78624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_110
timestamp 1669390400
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_111
timestamp 1669390400
transform -1 0 78624 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_112
timestamp 1669390400
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_113
timestamp 1669390400
transform -1 0 78624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_114
timestamp 1669390400
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_115
timestamp 1669390400
transform -1 0 78624 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_116
timestamp 1669390400
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_117
timestamp 1669390400
transform -1 0 78624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_118
timestamp 1669390400
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_119
timestamp 1669390400
transform -1 0 78624 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_120
timestamp 1669390400
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_121
timestamp 1669390400
transform -1 0 78624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_122
timestamp 1669390400
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_123
timestamp 1669390400
transform -1 0 78624 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_124
timestamp 1669390400
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_125
timestamp 1669390400
transform -1 0 78624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_126
timestamp 1669390400
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_127
timestamp 1669390400
transform -1 0 78624 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_128
timestamp 1669390400
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_129
timestamp 1669390400
transform -1 0 78624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_130
timestamp 1669390400
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_131
timestamp 1669390400
transform -1 0 78624 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_132
timestamp 1669390400
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_133
timestamp 1669390400
transform -1 0 78624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_134
timestamp 1669390400
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_135
timestamp 1669390400
transform -1 0 78624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_136
timestamp 1669390400
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_137
timestamp 1669390400
transform -1 0 78624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_138
timestamp 1669390400
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_139
timestamp 1669390400
transform -1 0 78624 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_140
timestamp 1669390400
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_141
timestamp 1669390400
transform -1 0 78624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_142
timestamp 1669390400
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_143
timestamp 1669390400
transform -1 0 78624 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_144
timestamp 1669390400
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_145
timestamp 1669390400
transform -1 0 78624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_146
timestamp 1669390400
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_147
timestamp 1669390400
transform -1 0 78624 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_148
timestamp 1669390400
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_149
timestamp 1669390400
transform -1 0 78624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_150
timestamp 1669390400
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_151
timestamp 1669390400
transform -1 0 78624 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_152
timestamp 1669390400
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_153
timestamp 1669390400
transform -1 0 78624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_154
timestamp 1669390400
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_155
timestamp 1669390400
transform -1 0 78624 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_156
timestamp 1669390400
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_157
timestamp 1669390400
transform -1 0 78624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_158
timestamp 1669390400
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_159
timestamp 1669390400
transform -1 0 78624 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_160
timestamp 1669390400
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_161
timestamp 1669390400
transform -1 0 78624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_162
timestamp 1669390400
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_163
timestamp 1669390400
transform -1 0 78624 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_164
timestamp 1669390400
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_165
timestamp 1669390400
transform -1 0 78624 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_166
timestamp 1669390400
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_167
timestamp 1669390400
transform -1 0 78624 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_168
timestamp 1669390400
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_169
timestamp 1669390400
transform -1 0 78624 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_170
timestamp 1669390400
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_171
timestamp 1669390400
transform -1 0 78624 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_172
timestamp 1669390400
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_173
timestamp 1669390400
transform -1 0 78624 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_174
timestamp 1669390400
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_175
timestamp 1669390400
transform -1 0 78624 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_176
timestamp 1669390400
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_177
timestamp 1669390400
transform -1 0 78624 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_178
timestamp 1669390400
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_179
timestamp 1669390400
transform -1 0 78624 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_180
timestamp 1669390400
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_181
timestamp 1669390400
transform -1 0 78624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_182
timestamp 1669390400
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_183
timestamp 1669390400
transform -1 0 78624 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_184
timestamp 1669390400
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_185
timestamp 1669390400
transform -1 0 78624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_186
timestamp 1669390400
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_187
timestamp 1669390400
transform -1 0 78624 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1669390400
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1669390400
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1669390400
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1669390400
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1669390400
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1669390400
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1669390400
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1669390400
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1669390400
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1669390400
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1669390400
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1669390400
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1669390400
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1669390400
transform 1 0 60144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1669390400
transform 1 0 64064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1669390400
transform 1 0 67984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1669390400
transform 1 0 71904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1669390400
transform 1 0 75824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1669390400
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1669390400
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1669390400
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1669390400
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1669390400
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1669390400
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1669390400
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1669390400
transform 1 0 64960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1669390400
transform 1 0 72912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1669390400
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1669390400
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1669390400
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1669390400
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1669390400
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1669390400
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1669390400
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1669390400
transform 1 0 60928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1669390400
transform 1 0 68880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1669390400
transform 1 0 76832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1669390400
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1669390400
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1669390400
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1669390400
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1669390400
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1669390400
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1669390400
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1669390400
transform 1 0 64960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1669390400
transform 1 0 72912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1669390400
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1669390400
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1669390400
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1669390400
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1669390400
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1669390400
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1669390400
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1669390400
transform 1 0 60928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1669390400
transform 1 0 68880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1669390400
transform 1 0 76832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1669390400
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1669390400
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1669390400
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1669390400
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1669390400
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1669390400
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1669390400
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1669390400
transform 1 0 64960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1669390400
transform 1 0 72912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1669390400
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1669390400
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1669390400
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1669390400
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1669390400
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1669390400
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1669390400
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1669390400
transform 1 0 60928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1669390400
transform 1 0 68880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1669390400
transform 1 0 76832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1669390400
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1669390400
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1669390400
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1669390400
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1669390400
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1669390400
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1669390400
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1669390400
transform 1 0 64960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1669390400
transform 1 0 72912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1669390400
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1669390400
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1669390400
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1669390400
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1669390400
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1669390400
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1669390400
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1669390400
transform 1 0 60928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1669390400
transform 1 0 68880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1669390400
transform 1 0 76832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1669390400
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1669390400
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1669390400
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1669390400
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1669390400
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1669390400
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1669390400
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1669390400
transform 1 0 64960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1669390400
transform 1 0 72912 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1669390400
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1669390400
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1669390400
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1669390400
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1669390400
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1669390400
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1669390400
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1669390400
transform 1 0 60928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1669390400
transform 1 0 68880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1669390400
transform 1 0 76832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1669390400
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1669390400
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1669390400
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1669390400
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1669390400
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1669390400
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1669390400
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1669390400
transform 1 0 64960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1669390400
transform 1 0 72912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1669390400
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1669390400
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1669390400
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1669390400
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1669390400
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1669390400
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1669390400
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1669390400
transform 1 0 60928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1669390400
transform 1 0 68880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1669390400
transform 1 0 76832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1669390400
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1669390400
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1669390400
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1669390400
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1669390400
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1669390400
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1669390400
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1669390400
transform 1 0 64960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1669390400
transform 1 0 72912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1669390400
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1669390400
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1669390400
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1669390400
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1669390400
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1669390400
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1669390400
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1669390400
transform 1 0 60928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1669390400
transform 1 0 68880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1669390400
transform 1 0 76832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1669390400
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1669390400
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1669390400
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1669390400
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1669390400
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1669390400
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1669390400
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1669390400
transform 1 0 64960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1669390400
transform 1 0 72912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1669390400
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1669390400
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1669390400
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1669390400
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1669390400
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1669390400
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1669390400
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1669390400
transform 1 0 60928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1669390400
transform 1 0 68880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1669390400
transform 1 0 76832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1669390400
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1669390400
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1669390400
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1669390400
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1669390400
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1669390400
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1669390400
transform 1 0 57008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1669390400
transform 1 0 64960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1669390400
transform 1 0 72912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1669390400
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1669390400
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1669390400
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1669390400
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1669390400
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1669390400
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1669390400
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1669390400
transform 1 0 60928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1669390400
transform 1 0 68880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1669390400
transform 1 0 76832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1669390400
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1669390400
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1669390400
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1669390400
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1669390400
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1669390400
transform 1 0 49056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1669390400
transform 1 0 57008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1669390400
transform 1 0 64960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1669390400
transform 1 0 72912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1669390400
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1669390400
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1669390400
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1669390400
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1669390400
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1669390400
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1669390400
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1669390400
transform 1 0 60928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1669390400
transform 1 0 68880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1669390400
transform 1 0 76832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1669390400
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1669390400
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1669390400
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1669390400
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1669390400
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1669390400
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1669390400
transform 1 0 57008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1669390400
transform 1 0 64960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1669390400
transform 1 0 72912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1669390400
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1669390400
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1669390400
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1669390400
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1669390400
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1669390400
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1669390400
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1669390400
transform 1 0 60928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1669390400
transform 1 0 68880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1669390400
transform 1 0 76832 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1669390400
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1669390400
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1669390400
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1669390400
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1669390400
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1669390400
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1669390400
transform 1 0 57008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1669390400
transform 1 0 64960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1669390400
transform 1 0 72912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1669390400
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1669390400
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1669390400
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1669390400
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1669390400
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1669390400
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1669390400
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1669390400
transform 1 0 60928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1669390400
transform 1 0 68880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1669390400
transform 1 0 76832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1669390400
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1669390400
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1669390400
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1669390400
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1669390400
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1669390400
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1669390400
transform 1 0 57008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1669390400
transform 1 0 64960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1669390400
transform 1 0 72912 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1669390400
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1669390400
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1669390400
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1669390400
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1669390400
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1669390400
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1669390400
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1669390400
transform 1 0 60928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1669390400
transform 1 0 68880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1669390400
transform 1 0 76832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1669390400
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1669390400
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1669390400
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1669390400
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1669390400
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1669390400
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1669390400
transform 1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1669390400
transform 1 0 64960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1669390400
transform 1 0 72912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1669390400
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1669390400
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1669390400
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1669390400
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1669390400
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1669390400
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1669390400
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1669390400
transform 1 0 60928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1669390400
transform 1 0 68880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1669390400
transform 1 0 76832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1669390400
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1669390400
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1669390400
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1669390400
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1669390400
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1669390400
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1669390400
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1669390400
transform 1 0 64960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1669390400
transform 1 0 72912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1669390400
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1669390400
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1669390400
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1669390400
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1669390400
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1669390400
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1669390400
transform 1 0 52976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1669390400
transform 1 0 60928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1669390400
transform 1 0 68880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1669390400
transform 1 0 76832 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1669390400
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1669390400
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1669390400
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1669390400
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1669390400
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1669390400
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1669390400
transform 1 0 57008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1669390400
transform 1 0 64960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1669390400
transform 1 0 72912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1669390400
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1669390400
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1669390400
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1669390400
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1669390400
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1669390400
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1669390400
transform 1 0 52976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1669390400
transform 1 0 60928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1669390400
transform 1 0 68880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1669390400
transform 1 0 76832 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1669390400
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1669390400
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_513
timestamp 1669390400
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_514
timestamp 1669390400
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_515
timestamp 1669390400
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_516
timestamp 1669390400
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_517
timestamp 1669390400
transform 1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_518
timestamp 1669390400
transform 1 0 64960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_519
timestamp 1669390400
transform 1 0 72912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_520
timestamp 1669390400
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_521
timestamp 1669390400
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_522
timestamp 1669390400
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_523
timestamp 1669390400
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_524
timestamp 1669390400
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_525
timestamp 1669390400
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_526
timestamp 1669390400
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_527
timestamp 1669390400
transform 1 0 60928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_528
timestamp 1669390400
transform 1 0 68880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_529
timestamp 1669390400
transform 1 0 76832 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_530
timestamp 1669390400
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_531
timestamp 1669390400
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_532
timestamp 1669390400
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_533
timestamp 1669390400
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_534
timestamp 1669390400
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_535
timestamp 1669390400
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_536
timestamp 1669390400
transform 1 0 57008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_537
timestamp 1669390400
transform 1 0 64960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_538
timestamp 1669390400
transform 1 0 72912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_539
timestamp 1669390400
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_540
timestamp 1669390400
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_541
timestamp 1669390400
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_542
timestamp 1669390400
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_543
timestamp 1669390400
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_544
timestamp 1669390400
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_545
timestamp 1669390400
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_546
timestamp 1669390400
transform 1 0 60928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_547
timestamp 1669390400
transform 1 0 68880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_548
timestamp 1669390400
transform 1 0 76832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_549
timestamp 1669390400
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_550
timestamp 1669390400
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_551
timestamp 1669390400
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_552
timestamp 1669390400
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_553
timestamp 1669390400
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_554
timestamp 1669390400
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_555
timestamp 1669390400
transform 1 0 57008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_556
timestamp 1669390400
transform 1 0 64960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_557
timestamp 1669390400
transform 1 0 72912 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_558
timestamp 1669390400
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_559
timestamp 1669390400
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_560
timestamp 1669390400
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_561
timestamp 1669390400
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_562
timestamp 1669390400
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_563
timestamp 1669390400
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_564
timestamp 1669390400
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_565
timestamp 1669390400
transform 1 0 60928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_566
timestamp 1669390400
transform 1 0 68880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_567
timestamp 1669390400
transform 1 0 76832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_568
timestamp 1669390400
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_569
timestamp 1669390400
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_570
timestamp 1669390400
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_571
timestamp 1669390400
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_572
timestamp 1669390400
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_573
timestamp 1669390400
transform 1 0 49056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_574
timestamp 1669390400
transform 1 0 57008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_575
timestamp 1669390400
transform 1 0 64960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_576
timestamp 1669390400
transform 1 0 72912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_577
timestamp 1669390400
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_578
timestamp 1669390400
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_579
timestamp 1669390400
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_580
timestamp 1669390400
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_581
timestamp 1669390400
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_582
timestamp 1669390400
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_583
timestamp 1669390400
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_584
timestamp 1669390400
transform 1 0 60928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_585
timestamp 1669390400
transform 1 0 68880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_586
timestamp 1669390400
transform 1 0 76832 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_587
timestamp 1669390400
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_588
timestamp 1669390400
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_589
timestamp 1669390400
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_590
timestamp 1669390400
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_591
timestamp 1669390400
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_592
timestamp 1669390400
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_593
timestamp 1669390400
transform 1 0 57008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_594
timestamp 1669390400
transform 1 0 64960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_595
timestamp 1669390400
transform 1 0 72912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_596
timestamp 1669390400
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_597
timestamp 1669390400
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_598
timestamp 1669390400
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_599
timestamp 1669390400
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_600
timestamp 1669390400
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_601
timestamp 1669390400
transform 1 0 45024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_602
timestamp 1669390400
transform 1 0 52976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_603
timestamp 1669390400
transform 1 0 60928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_604
timestamp 1669390400
transform 1 0 68880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_605
timestamp 1669390400
transform 1 0 76832 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_606
timestamp 1669390400
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_607
timestamp 1669390400
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_608
timestamp 1669390400
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_609
timestamp 1669390400
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_610
timestamp 1669390400
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_611
timestamp 1669390400
transform 1 0 49056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_612
timestamp 1669390400
transform 1 0 57008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_613
timestamp 1669390400
transform 1 0 64960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_614
timestamp 1669390400
transform 1 0 72912 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_615
timestamp 1669390400
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_616
timestamp 1669390400
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_617
timestamp 1669390400
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_618
timestamp 1669390400
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_619
timestamp 1669390400
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_620
timestamp 1669390400
transform 1 0 45024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_621
timestamp 1669390400
transform 1 0 52976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_622
timestamp 1669390400
transform 1 0 60928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_623
timestamp 1669390400
transform 1 0 68880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_624
timestamp 1669390400
transform 1 0 76832 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_625
timestamp 1669390400
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_626
timestamp 1669390400
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_627
timestamp 1669390400
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_628
timestamp 1669390400
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_629
timestamp 1669390400
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_630
timestamp 1669390400
transform 1 0 49056 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_631
timestamp 1669390400
transform 1 0 57008 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_632
timestamp 1669390400
transform 1 0 64960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_633
timestamp 1669390400
transform 1 0 72912 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_634
timestamp 1669390400
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_635
timestamp 1669390400
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_636
timestamp 1669390400
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_637
timestamp 1669390400
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_638
timestamp 1669390400
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_639
timestamp 1669390400
transform 1 0 45024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_640
timestamp 1669390400
transform 1 0 52976 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_641
timestamp 1669390400
transform 1 0 60928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_642
timestamp 1669390400
transform 1 0 68880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_643
timestamp 1669390400
transform 1 0 76832 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_644
timestamp 1669390400
transform 1 0 9296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_645
timestamp 1669390400
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_646
timestamp 1669390400
transform 1 0 25200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_647
timestamp 1669390400
transform 1 0 33152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_648
timestamp 1669390400
transform 1 0 41104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_649
timestamp 1669390400
transform 1 0 49056 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_650
timestamp 1669390400
transform 1 0 57008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_651
timestamp 1669390400
transform 1 0 64960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_652
timestamp 1669390400
transform 1 0 72912 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_653
timestamp 1669390400
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_654
timestamp 1669390400
transform 1 0 13216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_655
timestamp 1669390400
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_656
timestamp 1669390400
transform 1 0 29120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_657
timestamp 1669390400
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_658
timestamp 1669390400
transform 1 0 45024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_659
timestamp 1669390400
transform 1 0 52976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_660
timestamp 1669390400
transform 1 0 60928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_661
timestamp 1669390400
transform 1 0 68880 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_662
timestamp 1669390400
transform 1 0 76832 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_663
timestamp 1669390400
transform 1 0 9296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_664
timestamp 1669390400
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_665
timestamp 1669390400
transform 1 0 25200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_666
timestamp 1669390400
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_667
timestamp 1669390400
transform 1 0 41104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_668
timestamp 1669390400
transform 1 0 49056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_669
timestamp 1669390400
transform 1 0 57008 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_670
timestamp 1669390400
transform 1 0 64960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_671
timestamp 1669390400
transform 1 0 72912 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_672
timestamp 1669390400
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_673
timestamp 1669390400
transform 1 0 13216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_674
timestamp 1669390400
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_675
timestamp 1669390400
transform 1 0 29120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_676
timestamp 1669390400
transform 1 0 37072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_677
timestamp 1669390400
transform 1 0 45024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_678
timestamp 1669390400
transform 1 0 52976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_679
timestamp 1669390400
transform 1 0 60928 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_680
timestamp 1669390400
transform 1 0 68880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_681
timestamp 1669390400
transform 1 0 76832 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_682
timestamp 1669390400
transform 1 0 9296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_683
timestamp 1669390400
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_684
timestamp 1669390400
transform 1 0 25200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_685
timestamp 1669390400
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_686
timestamp 1669390400
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_687
timestamp 1669390400
transform 1 0 49056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_688
timestamp 1669390400
transform 1 0 57008 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_689
timestamp 1669390400
transform 1 0 64960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_690
timestamp 1669390400
transform 1 0 72912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_691
timestamp 1669390400
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_692
timestamp 1669390400
transform 1 0 13216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_693
timestamp 1669390400
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_694
timestamp 1669390400
transform 1 0 29120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_695
timestamp 1669390400
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_696
timestamp 1669390400
transform 1 0 45024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_697
timestamp 1669390400
transform 1 0 52976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_698
timestamp 1669390400
transform 1 0 60928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_699
timestamp 1669390400
transform 1 0 68880 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_700
timestamp 1669390400
transform 1 0 76832 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_701
timestamp 1669390400
transform 1 0 9296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_702
timestamp 1669390400
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_703
timestamp 1669390400
transform 1 0 25200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_704
timestamp 1669390400
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_705
timestamp 1669390400
transform 1 0 41104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_706
timestamp 1669390400
transform 1 0 49056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_707
timestamp 1669390400
transform 1 0 57008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_708
timestamp 1669390400
transform 1 0 64960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_709
timestamp 1669390400
transform 1 0 72912 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_710
timestamp 1669390400
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_711
timestamp 1669390400
transform 1 0 13216 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_712
timestamp 1669390400
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_713
timestamp 1669390400
transform 1 0 29120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_714
timestamp 1669390400
transform 1 0 37072 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_715
timestamp 1669390400
transform 1 0 45024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_716
timestamp 1669390400
transform 1 0 52976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_717
timestamp 1669390400
transform 1 0 60928 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_718
timestamp 1669390400
transform 1 0 68880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_719
timestamp 1669390400
transform 1 0 76832 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_720
timestamp 1669390400
transform 1 0 9296 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_721
timestamp 1669390400
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_722
timestamp 1669390400
transform 1 0 25200 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_723
timestamp 1669390400
transform 1 0 33152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_724
timestamp 1669390400
transform 1 0 41104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_725
timestamp 1669390400
transform 1 0 49056 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_726
timestamp 1669390400
transform 1 0 57008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_727
timestamp 1669390400
transform 1 0 64960 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_728
timestamp 1669390400
transform 1 0 72912 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_729
timestamp 1669390400
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_730
timestamp 1669390400
transform 1 0 13216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_731
timestamp 1669390400
transform 1 0 21168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_732
timestamp 1669390400
transform 1 0 29120 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_733
timestamp 1669390400
transform 1 0 37072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_734
timestamp 1669390400
transform 1 0 45024 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_735
timestamp 1669390400
transform 1 0 52976 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_736
timestamp 1669390400
transform 1 0 60928 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_737
timestamp 1669390400
transform 1 0 68880 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_738
timestamp 1669390400
transform 1 0 76832 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_739
timestamp 1669390400
transform 1 0 9296 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_740
timestamp 1669390400
transform 1 0 17248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_741
timestamp 1669390400
transform 1 0 25200 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_742
timestamp 1669390400
transform 1 0 33152 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_743
timestamp 1669390400
transform 1 0 41104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_744
timestamp 1669390400
transform 1 0 49056 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_745
timestamp 1669390400
transform 1 0 57008 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_746
timestamp 1669390400
transform 1 0 64960 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_747
timestamp 1669390400
transform 1 0 72912 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_748
timestamp 1669390400
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_749
timestamp 1669390400
transform 1 0 13216 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_750
timestamp 1669390400
transform 1 0 21168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_751
timestamp 1669390400
transform 1 0 29120 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_752
timestamp 1669390400
transform 1 0 37072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_753
timestamp 1669390400
transform 1 0 45024 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_754
timestamp 1669390400
transform 1 0 52976 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_755
timestamp 1669390400
transform 1 0 60928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_756
timestamp 1669390400
transform 1 0 68880 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_757
timestamp 1669390400
transform 1 0 76832 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_758
timestamp 1669390400
transform 1 0 9296 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_759
timestamp 1669390400
transform 1 0 17248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_760
timestamp 1669390400
transform 1 0 25200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_761
timestamp 1669390400
transform 1 0 33152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_762
timestamp 1669390400
transform 1 0 41104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_763
timestamp 1669390400
transform 1 0 49056 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_764
timestamp 1669390400
transform 1 0 57008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_765
timestamp 1669390400
transform 1 0 64960 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_766
timestamp 1669390400
transform 1 0 72912 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_767
timestamp 1669390400
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_768
timestamp 1669390400
transform 1 0 13216 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_769
timestamp 1669390400
transform 1 0 21168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_770
timestamp 1669390400
transform 1 0 29120 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_771
timestamp 1669390400
transform 1 0 37072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_772
timestamp 1669390400
transform 1 0 45024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_773
timestamp 1669390400
transform 1 0 52976 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_774
timestamp 1669390400
transform 1 0 60928 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_775
timestamp 1669390400
transform 1 0 68880 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_776
timestamp 1669390400
transform 1 0 76832 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_777
timestamp 1669390400
transform 1 0 9296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_778
timestamp 1669390400
transform 1 0 17248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_779
timestamp 1669390400
transform 1 0 25200 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_780
timestamp 1669390400
transform 1 0 33152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_781
timestamp 1669390400
transform 1 0 41104 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_782
timestamp 1669390400
transform 1 0 49056 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_783
timestamp 1669390400
transform 1 0 57008 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_784
timestamp 1669390400
transform 1 0 64960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_785
timestamp 1669390400
transform 1 0 72912 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_786
timestamp 1669390400
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_787
timestamp 1669390400
transform 1 0 13216 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_788
timestamp 1669390400
transform 1 0 21168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_789
timestamp 1669390400
transform 1 0 29120 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_790
timestamp 1669390400
transform 1 0 37072 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_791
timestamp 1669390400
transform 1 0 45024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_792
timestamp 1669390400
transform 1 0 52976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_793
timestamp 1669390400
transform 1 0 60928 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_794
timestamp 1669390400
transform 1 0 68880 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_795
timestamp 1669390400
transform 1 0 76832 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_796
timestamp 1669390400
transform 1 0 9296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_797
timestamp 1669390400
transform 1 0 17248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_798
timestamp 1669390400
transform 1 0 25200 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_799
timestamp 1669390400
transform 1 0 33152 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_800
timestamp 1669390400
transform 1 0 41104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_801
timestamp 1669390400
transform 1 0 49056 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_802
timestamp 1669390400
transform 1 0 57008 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_803
timestamp 1669390400
transform 1 0 64960 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_804
timestamp 1669390400
transform 1 0 72912 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_805
timestamp 1669390400
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_806
timestamp 1669390400
transform 1 0 13216 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_807
timestamp 1669390400
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_808
timestamp 1669390400
transform 1 0 29120 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_809
timestamp 1669390400
transform 1 0 37072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_810
timestamp 1669390400
transform 1 0 45024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_811
timestamp 1669390400
transform 1 0 52976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_812
timestamp 1669390400
transform 1 0 60928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_813
timestamp 1669390400
transform 1 0 68880 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_814
timestamp 1669390400
transform 1 0 76832 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_815
timestamp 1669390400
transform 1 0 9296 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_816
timestamp 1669390400
transform 1 0 17248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_817
timestamp 1669390400
transform 1 0 25200 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_818
timestamp 1669390400
transform 1 0 33152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_819
timestamp 1669390400
transform 1 0 41104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_820
timestamp 1669390400
transform 1 0 49056 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_821
timestamp 1669390400
transform 1 0 57008 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_822
timestamp 1669390400
transform 1 0 64960 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_823
timestamp 1669390400
transform 1 0 72912 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_824
timestamp 1669390400
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_825
timestamp 1669390400
transform 1 0 13216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_826
timestamp 1669390400
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_827
timestamp 1669390400
transform 1 0 29120 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_828
timestamp 1669390400
transform 1 0 37072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_829
timestamp 1669390400
transform 1 0 45024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_830
timestamp 1669390400
transform 1 0 52976 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_831
timestamp 1669390400
transform 1 0 60928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_832
timestamp 1669390400
transform 1 0 68880 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_833
timestamp 1669390400
transform 1 0 76832 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_834
timestamp 1669390400
transform 1 0 9296 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_835
timestamp 1669390400
transform 1 0 17248 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_836
timestamp 1669390400
transform 1 0 25200 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_837
timestamp 1669390400
transform 1 0 33152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_838
timestamp 1669390400
transform 1 0 41104 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_839
timestamp 1669390400
transform 1 0 49056 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_840
timestamp 1669390400
transform 1 0 57008 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_841
timestamp 1669390400
transform 1 0 64960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_842
timestamp 1669390400
transform 1 0 72912 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_843
timestamp 1669390400
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_844
timestamp 1669390400
transform 1 0 13216 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_845
timestamp 1669390400
transform 1 0 21168 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_846
timestamp 1669390400
transform 1 0 29120 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_847
timestamp 1669390400
transform 1 0 37072 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_848
timestamp 1669390400
transform 1 0 45024 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_849
timestamp 1669390400
transform 1 0 52976 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_850
timestamp 1669390400
transform 1 0 60928 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_851
timestamp 1669390400
transform 1 0 68880 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_852
timestamp 1669390400
transform 1 0 76832 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_853
timestamp 1669390400
transform 1 0 9296 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_854
timestamp 1669390400
transform 1 0 17248 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_855
timestamp 1669390400
transform 1 0 25200 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_856
timestamp 1669390400
transform 1 0 33152 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_857
timestamp 1669390400
transform 1 0 41104 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_858
timestamp 1669390400
transform 1 0 49056 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_859
timestamp 1669390400
transform 1 0 57008 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_860
timestamp 1669390400
transform 1 0 64960 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_861
timestamp 1669390400
transform 1 0 72912 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_862
timestamp 1669390400
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_863
timestamp 1669390400
transform 1 0 13216 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_864
timestamp 1669390400
transform 1 0 21168 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_865
timestamp 1669390400
transform 1 0 29120 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_866
timestamp 1669390400
transform 1 0 37072 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_867
timestamp 1669390400
transform 1 0 45024 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_868
timestamp 1669390400
transform 1 0 52976 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_869
timestamp 1669390400
transform 1 0 60928 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_870
timestamp 1669390400
transform 1 0 68880 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_871
timestamp 1669390400
transform 1 0 76832 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_872
timestamp 1669390400
transform 1 0 9296 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_873
timestamp 1669390400
transform 1 0 17248 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_874
timestamp 1669390400
transform 1 0 25200 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_875
timestamp 1669390400
transform 1 0 33152 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_876
timestamp 1669390400
transform 1 0 41104 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_877
timestamp 1669390400
transform 1 0 49056 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_878
timestamp 1669390400
transform 1 0 57008 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_879
timestamp 1669390400
transform 1 0 64960 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_880
timestamp 1669390400
transform 1 0 72912 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_881
timestamp 1669390400
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_882
timestamp 1669390400
transform 1 0 13216 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_883
timestamp 1669390400
transform 1 0 21168 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_884
timestamp 1669390400
transform 1 0 29120 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_885
timestamp 1669390400
transform 1 0 37072 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_886
timestamp 1669390400
transform 1 0 45024 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_887
timestamp 1669390400
transform 1 0 52976 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_888
timestamp 1669390400
transform 1 0 60928 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_889
timestamp 1669390400
transform 1 0 68880 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_890
timestamp 1669390400
transform 1 0 76832 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_891
timestamp 1669390400
transform 1 0 9296 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_892
timestamp 1669390400
transform 1 0 17248 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_893
timestamp 1669390400
transform 1 0 25200 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_894
timestamp 1669390400
transform 1 0 33152 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_895
timestamp 1669390400
transform 1 0 41104 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_896
timestamp 1669390400
transform 1 0 49056 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_897
timestamp 1669390400
transform 1 0 57008 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_898
timestamp 1669390400
transform 1 0 64960 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_899
timestamp 1669390400
transform 1 0 72912 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_900
timestamp 1669390400
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_901
timestamp 1669390400
transform 1 0 13216 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_902
timestamp 1669390400
transform 1 0 21168 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_903
timestamp 1669390400
transform 1 0 29120 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_904
timestamp 1669390400
transform 1 0 37072 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_905
timestamp 1669390400
transform 1 0 45024 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_906
timestamp 1669390400
transform 1 0 52976 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_907
timestamp 1669390400
transform 1 0 60928 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_908
timestamp 1669390400
transform 1 0 68880 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_909
timestamp 1669390400
transform 1 0 76832 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_910
timestamp 1669390400
transform 1 0 9296 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_911
timestamp 1669390400
transform 1 0 17248 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_912
timestamp 1669390400
transform 1 0 25200 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_913
timestamp 1669390400
transform 1 0 33152 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_914
timestamp 1669390400
transform 1 0 41104 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_915
timestamp 1669390400
transform 1 0 49056 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_916
timestamp 1669390400
transform 1 0 57008 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_917
timestamp 1669390400
transform 1 0 64960 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_918
timestamp 1669390400
transform 1 0 72912 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_919
timestamp 1669390400
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_920
timestamp 1669390400
transform 1 0 13216 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_921
timestamp 1669390400
transform 1 0 21168 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_922
timestamp 1669390400
transform 1 0 29120 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_923
timestamp 1669390400
transform 1 0 37072 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_924
timestamp 1669390400
transform 1 0 45024 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_925
timestamp 1669390400
transform 1 0 52976 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_926
timestamp 1669390400
transform 1 0 60928 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_927
timestamp 1669390400
transform 1 0 68880 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_928
timestamp 1669390400
transform 1 0 76832 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_929
timestamp 1669390400
transform 1 0 9296 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_930
timestamp 1669390400
transform 1 0 17248 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_931
timestamp 1669390400
transform 1 0 25200 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_932
timestamp 1669390400
transform 1 0 33152 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_933
timestamp 1669390400
transform 1 0 41104 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_934
timestamp 1669390400
transform 1 0 49056 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_935
timestamp 1669390400
transform 1 0 57008 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_936
timestamp 1669390400
transform 1 0 64960 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_937
timestamp 1669390400
transform 1 0 72912 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_938
timestamp 1669390400
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_939
timestamp 1669390400
transform 1 0 13216 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_940
timestamp 1669390400
transform 1 0 21168 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_941
timestamp 1669390400
transform 1 0 29120 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_942
timestamp 1669390400
transform 1 0 37072 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_943
timestamp 1669390400
transform 1 0 45024 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_944
timestamp 1669390400
transform 1 0 52976 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_945
timestamp 1669390400
transform 1 0 60928 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_946
timestamp 1669390400
transform 1 0 68880 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_947
timestamp 1669390400
transform 1 0 76832 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_948
timestamp 1669390400
transform 1 0 9296 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_949
timestamp 1669390400
transform 1 0 17248 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_950
timestamp 1669390400
transform 1 0 25200 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_951
timestamp 1669390400
transform 1 0 33152 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_952
timestamp 1669390400
transform 1 0 41104 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_953
timestamp 1669390400
transform 1 0 49056 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_954
timestamp 1669390400
transform 1 0 57008 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_955
timestamp 1669390400
transform 1 0 64960 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_956
timestamp 1669390400
transform 1 0 72912 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_957
timestamp 1669390400
transform 1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_958
timestamp 1669390400
transform 1 0 13216 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_959
timestamp 1669390400
transform 1 0 21168 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_960
timestamp 1669390400
transform 1 0 29120 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_961
timestamp 1669390400
transform 1 0 37072 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_962
timestamp 1669390400
transform 1 0 45024 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_963
timestamp 1669390400
transform 1 0 52976 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_964
timestamp 1669390400
transform 1 0 60928 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_965
timestamp 1669390400
transform 1 0 68880 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_966
timestamp 1669390400
transform 1 0 76832 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_967
timestamp 1669390400
transform 1 0 9296 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_968
timestamp 1669390400
transform 1 0 17248 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_969
timestamp 1669390400
transform 1 0 25200 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_970
timestamp 1669390400
transform 1 0 33152 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_971
timestamp 1669390400
transform 1 0 41104 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_972
timestamp 1669390400
transform 1 0 49056 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_973
timestamp 1669390400
transform 1 0 57008 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_974
timestamp 1669390400
transform 1 0 64960 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_975
timestamp 1669390400
transform 1 0 72912 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_976
timestamp 1669390400
transform 1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_977
timestamp 1669390400
transform 1 0 13216 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_978
timestamp 1669390400
transform 1 0 21168 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_979
timestamp 1669390400
transform 1 0 29120 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_980
timestamp 1669390400
transform 1 0 37072 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_981
timestamp 1669390400
transform 1 0 45024 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_982
timestamp 1669390400
transform 1 0 52976 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_983
timestamp 1669390400
transform 1 0 60928 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_984
timestamp 1669390400
transform 1 0 68880 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_985
timestamp 1669390400
transform 1 0 76832 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_986
timestamp 1669390400
transform 1 0 9296 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_987
timestamp 1669390400
transform 1 0 17248 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_988
timestamp 1669390400
transform 1 0 25200 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_989
timestamp 1669390400
transform 1 0 33152 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_990
timestamp 1669390400
transform 1 0 41104 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_991
timestamp 1669390400
transform 1 0 49056 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_992
timestamp 1669390400
transform 1 0 57008 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_993
timestamp 1669390400
transform 1 0 64960 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_994
timestamp 1669390400
transform 1 0 72912 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_995
timestamp 1669390400
transform 1 0 5264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_996
timestamp 1669390400
transform 1 0 13216 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_997
timestamp 1669390400
transform 1 0 21168 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_998
timestamp 1669390400
transform 1 0 29120 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_999
timestamp 1669390400
transform 1 0 37072 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1000
timestamp 1669390400
transform 1 0 45024 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1001
timestamp 1669390400
transform 1 0 52976 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1002
timestamp 1669390400
transform 1 0 60928 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1003
timestamp 1669390400
transform 1 0 68880 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1004
timestamp 1669390400
transform 1 0 76832 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1005
timestamp 1669390400
transform 1 0 9296 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1006
timestamp 1669390400
transform 1 0 17248 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1007
timestamp 1669390400
transform 1 0 25200 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1008
timestamp 1669390400
transform 1 0 33152 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1009
timestamp 1669390400
transform 1 0 41104 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1010
timestamp 1669390400
transform 1 0 49056 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1011
timestamp 1669390400
transform 1 0 57008 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1012
timestamp 1669390400
transform 1 0 64960 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1013
timestamp 1669390400
transform 1 0 72912 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1014
timestamp 1669390400
transform 1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1015
timestamp 1669390400
transform 1 0 13216 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1016
timestamp 1669390400
transform 1 0 21168 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1017
timestamp 1669390400
transform 1 0 29120 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1018
timestamp 1669390400
transform 1 0 37072 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1019
timestamp 1669390400
transform 1 0 45024 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1020
timestamp 1669390400
transform 1 0 52976 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1021
timestamp 1669390400
transform 1 0 60928 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1022
timestamp 1669390400
transform 1 0 68880 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1023
timestamp 1669390400
transform 1 0 76832 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1024
timestamp 1669390400
transform 1 0 9296 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1025
timestamp 1669390400
transform 1 0 17248 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1026
timestamp 1669390400
transform 1 0 25200 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1027
timestamp 1669390400
transform 1 0 33152 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1028
timestamp 1669390400
transform 1 0 41104 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1029
timestamp 1669390400
transform 1 0 49056 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1030
timestamp 1669390400
transform 1 0 57008 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1031
timestamp 1669390400
transform 1 0 64960 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1032
timestamp 1669390400
transform 1 0 72912 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1033
timestamp 1669390400
transform 1 0 5264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1034
timestamp 1669390400
transform 1 0 13216 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1035
timestamp 1669390400
transform 1 0 21168 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1036
timestamp 1669390400
transform 1 0 29120 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1037
timestamp 1669390400
transform 1 0 37072 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1038
timestamp 1669390400
transform 1 0 45024 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1039
timestamp 1669390400
transform 1 0 52976 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1040
timestamp 1669390400
transform 1 0 60928 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1041
timestamp 1669390400
transform 1 0 68880 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1042
timestamp 1669390400
transform 1 0 76832 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1043
timestamp 1669390400
transform 1 0 9296 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1044
timestamp 1669390400
transform 1 0 17248 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1045
timestamp 1669390400
transform 1 0 25200 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1046
timestamp 1669390400
transform 1 0 33152 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1047
timestamp 1669390400
transform 1 0 41104 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1048
timestamp 1669390400
transform 1 0 49056 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1049
timestamp 1669390400
transform 1 0 57008 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1050
timestamp 1669390400
transform 1 0 64960 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1051
timestamp 1669390400
transform 1 0 72912 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1052
timestamp 1669390400
transform 1 0 5264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1053
timestamp 1669390400
transform 1 0 13216 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1054
timestamp 1669390400
transform 1 0 21168 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1055
timestamp 1669390400
transform 1 0 29120 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1056
timestamp 1669390400
transform 1 0 37072 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1057
timestamp 1669390400
transform 1 0 45024 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1058
timestamp 1669390400
transform 1 0 52976 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1059
timestamp 1669390400
transform 1 0 60928 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1060
timestamp 1669390400
transform 1 0 68880 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1061
timestamp 1669390400
transform 1 0 76832 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1062
timestamp 1669390400
transform 1 0 9296 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1063
timestamp 1669390400
transform 1 0 17248 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1064
timestamp 1669390400
transform 1 0 25200 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1065
timestamp 1669390400
transform 1 0 33152 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1066
timestamp 1669390400
transform 1 0 41104 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1067
timestamp 1669390400
transform 1 0 49056 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1068
timestamp 1669390400
transform 1 0 57008 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1069
timestamp 1669390400
transform 1 0 64960 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1070
timestamp 1669390400
transform 1 0 72912 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1071
timestamp 1669390400
transform 1 0 5264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1072
timestamp 1669390400
transform 1 0 13216 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1073
timestamp 1669390400
transform 1 0 21168 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1074
timestamp 1669390400
transform 1 0 29120 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1075
timestamp 1669390400
transform 1 0 37072 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1076
timestamp 1669390400
transform 1 0 45024 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1077
timestamp 1669390400
transform 1 0 52976 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1078
timestamp 1669390400
transform 1 0 60928 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1079
timestamp 1669390400
transform 1 0 68880 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1080
timestamp 1669390400
transform 1 0 76832 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1081
timestamp 1669390400
transform 1 0 5264 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1082
timestamp 1669390400
transform 1 0 9184 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1083
timestamp 1669390400
transform 1 0 13104 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1084
timestamp 1669390400
transform 1 0 17024 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1085
timestamp 1669390400
transform 1 0 20944 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1086
timestamp 1669390400
transform 1 0 24864 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1087
timestamp 1669390400
transform 1 0 28784 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1088
timestamp 1669390400
transform 1 0 32704 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1089
timestamp 1669390400
transform 1 0 36624 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1090
timestamp 1669390400
transform 1 0 40544 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1091
timestamp 1669390400
transform 1 0 44464 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1092
timestamp 1669390400
transform 1 0 48384 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1093
timestamp 1669390400
transform 1 0 52304 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1094
timestamp 1669390400
transform 1 0 56224 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1095
timestamp 1669390400
transform 1 0 60144 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1096
timestamp 1669390400
transform 1 0 64064 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1097
timestamp 1669390400
transform 1 0 67984 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1098
timestamp 1669390400
transform 1 0 71904 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_1099
timestamp 1669390400
transform 1 0 75824 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _119_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 48720 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _120_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 44576 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _121_
timestamp 1669390400
transform 1 0 41664 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _122_
timestamp 1669390400
transform -1 0 46368 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _123_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 47040 0 -1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _124_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 45584 0 -1 73696
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _125_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 46704 0 1 72128
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _126_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 41888 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _127_
timestamp 1669390400
transform -1 0 47376 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _128_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 45584 0 1 73696
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _129_
timestamp 1669390400
transform -1 0 47152 0 -1 73696
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _130_
timestamp 1669390400
transform -1 0 43456 0 1 72128
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _131_
timestamp 1669390400
transform -1 0 39872 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _132_
timestamp 1669390400
transform 1 0 37520 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _133_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 45360 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _134_
timestamp 1669390400
transform -1 0 40208 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _135_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 38416 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _136_
timestamp 1669390400
transform -1 0 40544 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _137_
timestamp 1669390400
transform 1 0 37744 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _138_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 38192 0 1 72128
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _139_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 38416 0 -1 72128
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _140_
timestamp 1669390400
transform -1 0 44352 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _141_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 41888 0 -1 72128
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1669390400
transform -1 0 46256 0 -1 72128
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _143_
timestamp 1669390400
transform -1 0 45472 0 -1 72128
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _144_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 42448 0 -1 73696
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _145_
timestamp 1669390400
transform 1 0 43680 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _146_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 42560 0 1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _147_
timestamp 1669390400
transform -1 0 62496 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _148_
timestamp 1669390400
transform -1 0 56896 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _149_
timestamp 1669390400
transform -1 0 53536 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _150_
timestamp 1669390400
transform -1 0 60928 0 -1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _151_
timestamp 1669390400
transform -1 0 60144 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _152_
timestamp 1669390400
transform -1 0 56560 0 1 73696
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _153_
timestamp 1669390400
transform -1 0 52752 0 1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _154_
timestamp 1669390400
transform -1 0 52416 0 -1 75264
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _155_
timestamp 1669390400
transform -1 0 48944 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _156_
timestamp 1669390400
transform -1 0 60480 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _157_
timestamp 1669390400
transform -1 0 60032 0 1 73696
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _158_
timestamp 1669390400
transform -1 0 59808 0 -1 73696
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _159_
timestamp 1669390400
transform -1 0 54656 0 1 72128
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _160_
timestamp 1669390400
transform -1 0 59584 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _161_
timestamp 1669390400
transform 1 0 54992 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _162_
timestamp 1669390400
transform 1 0 59248 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _163_
timestamp 1669390400
transform -1 0 58016 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _164_
timestamp 1669390400
transform 1 0 55888 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _165_
timestamp 1669390400
transform -1 0 61600 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _166_
timestamp 1669390400
transform 1 0 56896 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _167_
timestamp 1669390400
transform 1 0 56112 0 1 70560
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _168_
timestamp 1669390400
transform 1 0 56336 0 1 72128
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _169_
timestamp 1669390400
transform -1 0 54656 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _170_
timestamp 1669390400
transform -1 0 54096 0 -1 73696
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _171_
timestamp 1669390400
transform 1 0 51408 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _172_
timestamp 1669390400
transform -1 0 51296 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _173_
timestamp 1669390400
transform 1 0 49504 0 -1 73696
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _174_
timestamp 1669390400
transform 1 0 49728 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _175_
timestamp 1669390400
transform -1 0 50736 0 1 73696
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _176_
timestamp 1669390400
transform 1 0 30912 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _177_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 50960 0 1 73696
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _178_
timestamp 1669390400
transform 1 0 43904 0 -1 75264
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _179_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 42896 0 -1 76832
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _180_
timestamp 1669390400
transform -1 0 35392 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _181_
timestamp 1669390400
transform -1 0 34720 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _182_
timestamp 1669390400
transform 1 0 36960 0 -1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _183_
timestamp 1669390400
transform 1 0 41440 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _184_
timestamp 1669390400
transform -1 0 46032 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _185_
timestamp 1669390400
transform -1 0 40096 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _186_
timestamp 1669390400
transform -1 0 40880 0 1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _187_
timestamp 1669390400
transform -1 0 61824 0 1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _188_
timestamp 1669390400
transform -1 0 57456 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _189_
timestamp 1669390400
transform -1 0 58352 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _190_
timestamp 1669390400
transform 1 0 55104 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _191_
timestamp 1669390400
transform -1 0 54544 0 1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _192_
timestamp 1669390400
transform 1 0 30016 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _193_
timestamp 1669390400
transform -1 0 30576 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _194_
timestamp 1669390400
transform -1 0 29008 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _195_
timestamp 1669390400
transform -1 0 31696 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _196_
timestamp 1669390400
transform 1 0 29792 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _197_
timestamp 1669390400
transform -1 0 31696 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _198_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 30688 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _199_
timestamp 1669390400
transform -1 0 39424 0 -1 73696
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _200_
timestamp 1669390400
transform 1 0 38752 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _201_
timestamp 1669390400
transform -1 0 37968 0 1 72128
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _202_
timestamp 1669390400
transform 1 0 36400 0 1 72128
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _203_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 40992 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _204_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 36176 0 -1 73696
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _205_
timestamp 1669390400
transform 1 0 57456 0 -1 72128
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _206_
timestamp 1669390400
transform 1 0 55888 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _207_
timestamp 1669390400
transform 1 0 57792 0 1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _208_
timestamp 1669390400
transform -1 0 60816 0 1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _209_
timestamp 1669390400
transform -1 0 59248 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _210_
timestamp 1669390400
transform 1 0 57344 0 -1 75264
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _211_
timestamp 1669390400
transform 1 0 32704 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _212_
timestamp 1669390400
transform -1 0 34160 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _213_
timestamp 1669390400
transform -1 0 33040 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _214_
timestamp 1669390400
transform 1 0 31920 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _215_
timestamp 1669390400
transform -1 0 32480 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _216_
timestamp 1669390400
transform -1 0 34608 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _217_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 40544 0 1 70560
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _218_
timestamp 1669390400
transform 1 0 38304 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _219_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 42560 0 -1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _220_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 44688 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _221_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 41664 0 1 73696
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _222_
timestamp 1669390400
transform 1 0 51408 0 1 72128
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _223_
timestamp 1669390400
transform -1 0 55552 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _224_
timestamp 1669390400
transform 1 0 53760 0 -1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _225_
timestamp 1669390400
transform -1 0 55216 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _226_
timestamp 1669390400
transform 1 0 53312 0 1 73696
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _227_
timestamp 1669390400
transform 1 0 34384 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _228_
timestamp 1669390400
transform 1 0 35168 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _229_
timestamp 1669390400
transform 1 0 34048 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _230_
timestamp 1669390400
transform 1 0 42336 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _231_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 44912 0 1 70560
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _232_
timestamp 1669390400
transform -1 0 42000 0 -1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _233_
timestamp 1669390400
transform 1 0 40432 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _234_
timestamp 1669390400
transform 1 0 36400 0 1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _235_
timestamp 1669390400
transform 1 0 36288 0 -1 75264
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _236_
timestamp 1669390400
transform 1 0 52304 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _237_
timestamp 1669390400
transform -1 0 52080 0 -1 72128
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _238_
timestamp 1669390400
transform -1 0 51296 0 -1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _239_
timestamp 1669390400
transform -1 0 51184 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _240_
timestamp 1669390400
transform -1 0 49280 0 -1 76832
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _241_
timestamp 1669390400
transform 1 0 47264 0 -1 75264
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _242_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 49504 0 -1 76832
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _243_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 50512 0 -1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _244_
timestamp 1669390400
transform -1 0 40992 0 -1 73696
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _245_
timestamp 1669390400
transform -1 0 38528 0 1 73696
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _246_
timestamp 1669390400
transform -1 0 36960 0 1 75264
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _247_
timestamp 1669390400
transform -1 0 34944 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _248_
timestamp 1669390400
transform -1 0 29568 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _249_
timestamp 1669390400
transform 1 0 30240 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _250_
timestamp 1669390400
transform -1 0 36064 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _251_
timestamp 1669390400
transform -1 0 35728 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _252_
timestamp 1669390400
transform 1 0 36848 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input1 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1680 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input2
timestamp 1669390400
transform 1 0 38640 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input3
timestamp 1669390400
transform -1 0 42672 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1669390400
transform -1 0 45472 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input5
timestamp 1669390400
transform -1 0 47264 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input6 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 49504 0 1 75264
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1669390400
transform -1 0 48272 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input8
timestamp 1669390400
transform -1 0 55440 0 -1 76832
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input9
timestamp 1669390400
transform -1 0 52192 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input10
timestamp 1669390400
transform 1 0 54768 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input11
timestamp 1669390400
transform -1 0 58576 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1669390400
transform -1 0 59472 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input13
timestamp 1669390400
transform -1 0 61488 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input14
timestamp 1669390400
transform -1 0 65632 0 1 75264
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input15
timestamp 1669390400
transform -1 0 67648 0 -1 76832
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input16
timestamp 1669390400
transform -1 0 71120 0 -1 76832
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input17
timestamp 1669390400
transform -1 0 69888 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input18
timestamp 1669390400
transform -1 0 73696 0 1 75264
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1669390400
transform -1 0 73584 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input20
timestamp 1669390400
transform -1 0 76720 0 1 75264
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyd_1  input21 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 78288 0 -1 75264
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_37 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 55776 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_38
timestamp 1669390400
transform -1 0 55664 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_39
timestamp 1669390400
transform -1 0 57008 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_40
timestamp 1669390400
transform -1 0 57680 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_41
timestamp 1669390400
transform -1 0 58352 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_42
timestamp 1669390400
transform -1 0 59024 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_43
timestamp 1669390400
transform -1 0 59696 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_44
timestamp 1669390400
transform -1 0 59696 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_45
timestamp 1669390400
transform -1 0 60928 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_46
timestamp 1669390400
transform -1 0 61600 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_47
timestamp 1669390400
transform -1 0 62272 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_48
timestamp 1669390400
transform -1 0 62944 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_49
timestamp 1669390400
transform -1 0 63616 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_50
timestamp 1669390400
transform -1 0 63728 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_51
timestamp 1669390400
transform -1 0 64848 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_52
timestamp 1669390400
transform -1 0 65520 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_53
timestamp 1669390400
transform -1 0 66192 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_54
timestamp 1669390400
transform -1 0 66864 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_55
timestamp 1669390400
transform -1 0 67536 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_56
timestamp 1669390400
transform -1 0 68768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_57
timestamp 1669390400
transform -1 0 69440 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_58
timestamp 1669390400
transform -1 0 70112 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_59
timestamp 1669390400
transform -1 0 70784 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_60
timestamp 1669390400
transform -1 0 71456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_61
timestamp 1669390400
transform -1 0 71120 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_62
timestamp 1669390400
transform -1 0 72688 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_63
timestamp 1669390400
transform -1 0 73360 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_64
timestamp 1669390400
transform -1 0 74032 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_65
timestamp 1669390400
transform -1 0 7280 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_66
timestamp 1669390400
transform -1 0 8400 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_67
timestamp 1669390400
transform 1 0 8624 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_68
timestamp 1669390400
transform -1 0 10304 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_69
timestamp 1669390400
transform 1 0 10528 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_70
timestamp 1669390400
transform 1 0 11200 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_71
timestamp 1669390400
transform 1 0 11872 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_72
timestamp 1669390400
transform 1 0 12544 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_73
timestamp 1669390400
transform -1 0 14224 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_74
timestamp 1669390400
transform 1 0 13776 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_75
timestamp 1669390400
transform 1 0 14448 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_76
timestamp 1669390400
transform 1 0 15120 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_77
timestamp 1669390400
transform 1 0 15792 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_78
timestamp 1669390400
transform 1 0 16464 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_79
timestamp 1669390400
transform -1 0 18256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_80
timestamp 1669390400
transform 1 0 17696 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_81
timestamp 1669390400
transform 1 0 18368 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_82
timestamp 1669390400
transform 1 0 19040 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_83
timestamp 1669390400
transform 1 0 19712 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_84
timestamp 1669390400
transform 1 0 20384 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_85
timestamp 1669390400
transform -1 0 22064 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_86
timestamp 1669390400
transform -1 0 22736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_87
timestamp 1669390400
transform -1 0 23408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_88
timestamp 1669390400
transform -1 0 24080 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_89
timestamp 1669390400
transform -1 0 24976 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_90
timestamp 1669390400
transform 1 0 24304 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_91
timestamp 1669390400
transform 1 0 25536 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_92
timestamp 1669390400
transform 1 0 26208 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_93
timestamp 1669390400
transform 1 0 26880 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_94
timestamp 1669390400
transform 1 0 27552 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_95
timestamp 1669390400
transform 1 0 28224 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_96
timestamp 1669390400
transform -1 0 29680 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_97
timestamp 1669390400
transform 1 0 29456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_98
timestamp 1669390400
transform -1 0 4144 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_99
timestamp 1669390400
transform 1 0 4704 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_100
timestamp 1669390400
transform -1 0 7504 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_101
timestamp 1669390400
transform 1 0 8624 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_102
timestamp 1669390400
transform 1 0 10752 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_103
timestamp 1669390400
transform -1 0 14000 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_104
timestamp 1669390400
transform -1 0 15568 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_105
timestamp 1669390400
transform -1 0 17584 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_106
timestamp 1669390400
transform -1 0 19600 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_107
timestamp 1669390400
transform -1 0 21952 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_108
timestamp 1669390400
transform -1 0 23632 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_109
timestamp 1669390400
transform -1 0 25648 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_110
timestamp 1669390400
transform -1 0 27440 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_111
timestamp 1669390400
transform 1 0 27664 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_112
timestamp 1669390400
transform -1 0 32368 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_113
timestamp 1669390400
transform 1 0 29232 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_114
timestamp 1669390400
transform -1 0 35728 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_115
timestamp 1669390400
transform 1 0 35728 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_116
timestamp 1669390400
transform 1 0 38752 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_117
timestamp 1669390400
transform -1 0 41888 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_118
timestamp 1669390400
transform -1 0 48048 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_119
timestamp 1669390400
transform -1 0 49392 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_120
timestamp 1669390400
transform -1 0 48048 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_121
timestamp 1669390400
transform -1 0 56112 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_122
timestamp 1669390400
transform -1 0 51856 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_123
timestamp 1669390400
transform -1 0 53872 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_124
timestamp 1669390400
transform -1 0 62160 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_125
timestamp 1669390400
transform -1 0 63504 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_126
timestamp 1669390400
transform -1 0 61712 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_127
timestamp 1669390400
transform -1 0 62944 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_128
timestamp 1669390400
transform -1 0 64288 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_129
timestamp 1669390400
transform -1 0 66976 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_130
timestamp 1669390400
transform -1 0 68320 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_131
timestamp 1669390400
transform -1 0 70560 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_132
timestamp 1669390400
transform -1 0 72688 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_133
timestamp 1669390400
transform -1 0 74928 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_134
timestamp 1669390400
transform -1 0 76608 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_135
timestamp 1669390400
transform -1 0 78064 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_136
timestamp 1669390400
transform -1 0 6160 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_137
timestamp 1669390400
transform -1 0 8176 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_138
timestamp 1669390400
transform -1 0 10192 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_139
timestamp 1669390400
transform 1 0 35504 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_140
timestamp 1669390400
transform -1 0 47376 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_141
timestamp 1669390400
transform -1 0 47824 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_142
timestamp 1669390400
transform -1 0 46928 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_143
timestamp 1669390400
transform -1 0 48720 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_144
timestamp 1669390400
transform 1 0 49056 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_145
timestamp 1669390400
transform -1 0 52528 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_146
timestamp 1669390400
transform -1 0 60816 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_147
timestamp 1669390400
transform -1 0 62832 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_148
timestamp 1669390400
transform -1 0 62272 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_149
timestamp 1669390400
transform -1 0 61152 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_150
timestamp 1669390400
transform -1 0 63616 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_151
timestamp 1669390400
transform -1 0 66304 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_152
timestamp 1669390400
transform -1 0 67648 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_153
timestamp 1669390400
transform -1 0 68656 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_154
timestamp 1669390400
transform -1 0 71792 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_155
timestamp 1669390400
transform -1 0 74256 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_156
timestamp 1669390400
transform -1 0 75600 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_157
timestamp 1669390400
transform -1 0 77280 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_158
timestamp 1669390400
transform 1 0 77840 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_159
timestamp 1669390400
transform -1 0 73696 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_160
timestamp 1669390400
transform -1 0 74704 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_161
timestamp 1669390400
transform -1 0 74368 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_162
timestamp 1669390400
transform -1 0 30576 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_163
timestamp 1669390400
transform -1 0 31248 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_164
timestamp 1669390400
transform -1 0 31920 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_165
timestamp 1669390400
transform -1 0 32816 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_166
timestamp 1669390400
transform 1 0 32144 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_167
timestamp 1669390400
transform 1 0 33376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_168
timestamp 1669390400
transform 1 0 34048 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_169
timestamp 1669390400
transform 1 0 34720 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_170
timestamp 1669390400
transform 1 0 35392 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_171
timestamp 1669390400
transform 1 0 36064 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_172
timestamp 1669390400
transform -1 0 37520 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_173
timestamp 1669390400
transform 1 0 37296 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_174
timestamp 1669390400
transform 1 0 37968 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_175
timestamp 1669390400
transform 1 0 38640 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_176
timestamp 1669390400
transform 1 0 39312 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_177
timestamp 1669390400
transform 1 0 39984 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_178
timestamp 1669390400
transform -1 0 41552 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_179
timestamp 1669390400
transform -1 0 42224 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_180
timestamp 1669390400
transform -1 0 42896 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_181
timestamp 1669390400
transform -1 0 43568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_182
timestamp 1669390400
transform -1 0 44240 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_183
timestamp 1669390400
transform -1 0 45248 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_184
timestamp 1669390400
transform -1 0 45920 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_185
timestamp 1669390400
transform -1 0 46592 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_186
timestamp 1669390400
transform -1 0 47264 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_187
timestamp 1669390400
transform -1 0 47936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_188
timestamp 1669390400
transform -1 0 49168 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_189
timestamp 1669390400
transform -1 0 49840 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_190
timestamp 1669390400
transform -1 0 50512 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_191
timestamp 1669390400
transform -1 0 51184 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_192
timestamp 1669390400
transform -1 0 51856 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_193
timestamp 1669390400
transform -1 0 51632 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_194
timestamp 1669390400
transform -1 0 53088 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_195
timestamp 1669390400
transform -1 0 53760 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_196
timestamp 1669390400
transform -1 0 54432 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_decap64_197
timestamp 1669390400
transform -1 0 55104 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output22 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 7168 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output23
timestamp 1669390400
transform -1 0 24752 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output24
timestamp 1669390400
transform -1 0 26880 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output25
timestamp 1669390400
transform -1 0 28672 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output26
timestamp 1669390400
transform -1 0 31472 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output27
timestamp 1669390400
transform 1 0 31920 0 1 75264
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output28
timestamp 1669390400
transform 1 0 33152 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output29
timestamp 1669390400
transform 1 0 34944 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output30
timestamp 1669390400
transform 1 0 37968 0 1 75264
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output31
timestamp 1669390400
transform -1 0 12992 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output32
timestamp 1669390400
transform -1 0 15120 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output33
timestamp 1669390400
transform -1 0 16912 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output34
timestamp 1669390400
transform -1 0 19040 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output35
timestamp 1669390400
transform -1 0 20832 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output36
timestamp 1669390400
transform -1 0 22960 0 -1 76832
box -86 -86 1654 870
<< labels >>
flabel metal2 s 1568 79200 1680 80000 0 FreeSans 448 90 0 0 io_active
port 0 nsew signal input
flabel metal2 s 2240 79200 2352 80000 0 FreeSans 448 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 22400 79200 22512 80000 0 FreeSans 448 90 0 0 io_in[10]
port 2 nsew signal input
flabel metal2 s 24416 79200 24528 80000 0 FreeSans 448 90 0 0 io_in[11]
port 3 nsew signal input
flabel metal2 s 26432 79200 26544 80000 0 FreeSans 448 90 0 0 io_in[12]
port 4 nsew signal input
flabel metal2 s 28448 79200 28560 80000 0 FreeSans 448 90 0 0 io_in[13]
port 5 nsew signal input
flabel metal2 s 30464 79200 30576 80000 0 FreeSans 448 90 0 0 io_in[14]
port 6 nsew signal input
flabel metal2 s 32480 79200 32592 80000 0 FreeSans 448 90 0 0 io_in[15]
port 7 nsew signal input
flabel metal2 s 34496 79200 34608 80000 0 FreeSans 448 90 0 0 io_in[16]
port 8 nsew signal input
flabel metal2 s 36512 79200 36624 80000 0 FreeSans 448 90 0 0 io_in[17]
port 9 nsew signal input
flabel metal2 s 38528 79200 38640 80000 0 FreeSans 448 90 0 0 io_in[18]
port 10 nsew signal input
flabel metal2 s 40544 79200 40656 80000 0 FreeSans 448 90 0 0 io_in[19]
port 11 nsew signal input
flabel metal2 s 4256 79200 4368 80000 0 FreeSans 448 90 0 0 io_in[1]
port 12 nsew signal input
flabel metal2 s 42560 79200 42672 80000 0 FreeSans 448 90 0 0 io_in[20]
port 13 nsew signal input
flabel metal2 s 44576 79200 44688 80000 0 FreeSans 448 90 0 0 io_in[21]
port 14 nsew signal input
flabel metal2 s 46592 79200 46704 80000 0 FreeSans 448 90 0 0 io_in[22]
port 15 nsew signal input
flabel metal2 s 48608 79200 48720 80000 0 FreeSans 448 90 0 0 io_in[23]
port 16 nsew signal input
flabel metal2 s 50624 79200 50736 80000 0 FreeSans 448 90 0 0 io_in[24]
port 17 nsew signal input
flabel metal2 s 52640 79200 52752 80000 0 FreeSans 448 90 0 0 io_in[25]
port 18 nsew signal input
flabel metal2 s 54656 79200 54768 80000 0 FreeSans 448 90 0 0 io_in[26]
port 19 nsew signal input
flabel metal2 s 56672 79200 56784 80000 0 FreeSans 448 90 0 0 io_in[27]
port 20 nsew signal input
flabel metal2 s 58688 79200 58800 80000 0 FreeSans 448 90 0 0 io_in[28]
port 21 nsew signal input
flabel metal2 s 60704 79200 60816 80000 0 FreeSans 448 90 0 0 io_in[29]
port 22 nsew signal input
flabel metal2 s 6272 79200 6384 80000 0 FreeSans 448 90 0 0 io_in[2]
port 23 nsew signal input
flabel metal2 s 62720 79200 62832 80000 0 FreeSans 448 90 0 0 io_in[30]
port 24 nsew signal input
flabel metal2 s 64736 79200 64848 80000 0 FreeSans 448 90 0 0 io_in[31]
port 25 nsew signal input
flabel metal2 s 66752 79200 66864 80000 0 FreeSans 448 90 0 0 io_in[32]
port 26 nsew signal input
flabel metal2 s 68768 79200 68880 80000 0 FreeSans 448 90 0 0 io_in[33]
port 27 nsew signal input
flabel metal2 s 70784 79200 70896 80000 0 FreeSans 448 90 0 0 io_in[34]
port 28 nsew signal input
flabel metal2 s 72800 79200 72912 80000 0 FreeSans 448 90 0 0 io_in[35]
port 29 nsew signal input
flabel metal2 s 74816 79200 74928 80000 0 FreeSans 448 90 0 0 io_in[36]
port 30 nsew signal input
flabel metal2 s 76832 79200 76944 80000 0 FreeSans 448 90 0 0 io_in[37]
port 31 nsew signal input
flabel metal2 s 8288 79200 8400 80000 0 FreeSans 448 90 0 0 io_in[3]
port 32 nsew signal input
flabel metal2 s 10304 79200 10416 80000 0 FreeSans 448 90 0 0 io_in[4]
port 33 nsew signal input
flabel metal2 s 12320 79200 12432 80000 0 FreeSans 448 90 0 0 io_in[5]
port 34 nsew signal input
flabel metal2 s 14336 79200 14448 80000 0 FreeSans 448 90 0 0 io_in[6]
port 35 nsew signal input
flabel metal2 s 16352 79200 16464 80000 0 FreeSans 448 90 0 0 io_in[7]
port 36 nsew signal input
flabel metal2 s 18368 79200 18480 80000 0 FreeSans 448 90 0 0 io_in[8]
port 37 nsew signal input
flabel metal2 s 20384 79200 20496 80000 0 FreeSans 448 90 0 0 io_in[9]
port 38 nsew signal input
flabel metal2 s 2912 79200 3024 80000 0 FreeSans 448 90 0 0 io_oeb[0]
port 39 nsew signal tristate
flabel metal2 s 23072 79200 23184 80000 0 FreeSans 448 90 0 0 io_oeb[10]
port 40 nsew signal tristate
flabel metal2 s 25088 79200 25200 80000 0 FreeSans 448 90 0 0 io_oeb[11]
port 41 nsew signal tristate
flabel metal2 s 27104 79200 27216 80000 0 FreeSans 448 90 0 0 io_oeb[12]
port 42 nsew signal tristate
flabel metal2 s 29120 79200 29232 80000 0 FreeSans 448 90 0 0 io_oeb[13]
port 43 nsew signal tristate
flabel metal2 s 31136 79200 31248 80000 0 FreeSans 448 90 0 0 io_oeb[14]
port 44 nsew signal tristate
flabel metal2 s 33152 79200 33264 80000 0 FreeSans 448 90 0 0 io_oeb[15]
port 45 nsew signal tristate
flabel metal2 s 35168 79200 35280 80000 0 FreeSans 448 90 0 0 io_oeb[16]
port 46 nsew signal tristate
flabel metal2 s 37184 79200 37296 80000 0 FreeSans 448 90 0 0 io_oeb[17]
port 47 nsew signal tristate
flabel metal2 s 39200 79200 39312 80000 0 FreeSans 448 90 0 0 io_oeb[18]
port 48 nsew signal tristate
flabel metal2 s 41216 79200 41328 80000 0 FreeSans 448 90 0 0 io_oeb[19]
port 49 nsew signal tristate
flabel metal2 s 4928 79200 5040 80000 0 FreeSans 448 90 0 0 io_oeb[1]
port 50 nsew signal tristate
flabel metal2 s 43232 79200 43344 80000 0 FreeSans 448 90 0 0 io_oeb[20]
port 51 nsew signal tristate
flabel metal2 s 45248 79200 45360 80000 0 FreeSans 448 90 0 0 io_oeb[21]
port 52 nsew signal tristate
flabel metal2 s 47264 79200 47376 80000 0 FreeSans 448 90 0 0 io_oeb[22]
port 53 nsew signal tristate
flabel metal2 s 49280 79200 49392 80000 0 FreeSans 448 90 0 0 io_oeb[23]
port 54 nsew signal tristate
flabel metal2 s 51296 79200 51408 80000 0 FreeSans 448 90 0 0 io_oeb[24]
port 55 nsew signal tristate
flabel metal2 s 53312 79200 53424 80000 0 FreeSans 448 90 0 0 io_oeb[25]
port 56 nsew signal tristate
flabel metal2 s 55328 79200 55440 80000 0 FreeSans 448 90 0 0 io_oeb[26]
port 57 nsew signal tristate
flabel metal2 s 57344 79200 57456 80000 0 FreeSans 448 90 0 0 io_oeb[27]
port 58 nsew signal tristate
flabel metal2 s 59360 79200 59472 80000 0 FreeSans 448 90 0 0 io_oeb[28]
port 59 nsew signal tristate
flabel metal2 s 61376 79200 61488 80000 0 FreeSans 448 90 0 0 io_oeb[29]
port 60 nsew signal tristate
flabel metal2 s 6944 79200 7056 80000 0 FreeSans 448 90 0 0 io_oeb[2]
port 61 nsew signal tristate
flabel metal2 s 63392 79200 63504 80000 0 FreeSans 448 90 0 0 io_oeb[30]
port 62 nsew signal tristate
flabel metal2 s 65408 79200 65520 80000 0 FreeSans 448 90 0 0 io_oeb[31]
port 63 nsew signal tristate
flabel metal2 s 67424 79200 67536 80000 0 FreeSans 448 90 0 0 io_oeb[32]
port 64 nsew signal tristate
flabel metal2 s 69440 79200 69552 80000 0 FreeSans 448 90 0 0 io_oeb[33]
port 65 nsew signal tristate
flabel metal2 s 71456 79200 71568 80000 0 FreeSans 448 90 0 0 io_oeb[34]
port 66 nsew signal tristate
flabel metal2 s 73472 79200 73584 80000 0 FreeSans 448 90 0 0 io_oeb[35]
port 67 nsew signal tristate
flabel metal2 s 75488 79200 75600 80000 0 FreeSans 448 90 0 0 io_oeb[36]
port 68 nsew signal tristate
flabel metal2 s 77504 79200 77616 80000 0 FreeSans 448 90 0 0 io_oeb[37]
port 69 nsew signal tristate
flabel metal2 s 8960 79200 9072 80000 0 FreeSans 448 90 0 0 io_oeb[3]
port 70 nsew signal tristate
flabel metal2 s 10976 79200 11088 80000 0 FreeSans 448 90 0 0 io_oeb[4]
port 71 nsew signal tristate
flabel metal2 s 12992 79200 13104 80000 0 FreeSans 448 90 0 0 io_oeb[5]
port 72 nsew signal tristate
flabel metal2 s 15008 79200 15120 80000 0 FreeSans 448 90 0 0 io_oeb[6]
port 73 nsew signal tristate
flabel metal2 s 17024 79200 17136 80000 0 FreeSans 448 90 0 0 io_oeb[7]
port 74 nsew signal tristate
flabel metal2 s 19040 79200 19152 80000 0 FreeSans 448 90 0 0 io_oeb[8]
port 75 nsew signal tristate
flabel metal2 s 21056 79200 21168 80000 0 FreeSans 448 90 0 0 io_oeb[9]
port 76 nsew signal tristate
flabel metal2 s 3584 79200 3696 80000 0 FreeSans 448 90 0 0 io_out[0]
port 77 nsew signal tristate
flabel metal2 s 23744 79200 23856 80000 0 FreeSans 448 90 0 0 io_out[10]
port 78 nsew signal tristate
flabel metal2 s 25760 79200 25872 80000 0 FreeSans 448 90 0 0 io_out[11]
port 79 nsew signal tristate
flabel metal2 s 27776 79200 27888 80000 0 FreeSans 448 90 0 0 io_out[12]
port 80 nsew signal tristate
flabel metal2 s 29792 79200 29904 80000 0 FreeSans 448 90 0 0 io_out[13]
port 81 nsew signal tristate
flabel metal2 s 31808 79200 31920 80000 0 FreeSans 448 90 0 0 io_out[14]
port 82 nsew signal tristate
flabel metal2 s 33824 79200 33936 80000 0 FreeSans 448 90 0 0 io_out[15]
port 83 nsew signal tristate
flabel metal2 s 35840 79200 35952 80000 0 FreeSans 448 90 0 0 io_out[16]
port 84 nsew signal tristate
flabel metal2 s 37856 79200 37968 80000 0 FreeSans 448 90 0 0 io_out[17]
port 85 nsew signal tristate
flabel metal2 s 39872 79200 39984 80000 0 FreeSans 448 90 0 0 io_out[18]
port 86 nsew signal tristate
flabel metal2 s 41888 79200 42000 80000 0 FreeSans 448 90 0 0 io_out[19]
port 87 nsew signal tristate
flabel metal2 s 5600 79200 5712 80000 0 FreeSans 448 90 0 0 io_out[1]
port 88 nsew signal tristate
flabel metal2 s 43904 79200 44016 80000 0 FreeSans 448 90 0 0 io_out[20]
port 89 nsew signal tristate
flabel metal2 s 45920 79200 46032 80000 0 FreeSans 448 90 0 0 io_out[21]
port 90 nsew signal tristate
flabel metal2 s 47936 79200 48048 80000 0 FreeSans 448 90 0 0 io_out[22]
port 91 nsew signal tristate
flabel metal2 s 49952 79200 50064 80000 0 FreeSans 448 90 0 0 io_out[23]
port 92 nsew signal tristate
flabel metal2 s 51968 79200 52080 80000 0 FreeSans 448 90 0 0 io_out[24]
port 93 nsew signal tristate
flabel metal2 s 53984 79200 54096 80000 0 FreeSans 448 90 0 0 io_out[25]
port 94 nsew signal tristate
flabel metal2 s 56000 79200 56112 80000 0 FreeSans 448 90 0 0 io_out[26]
port 95 nsew signal tristate
flabel metal2 s 58016 79200 58128 80000 0 FreeSans 448 90 0 0 io_out[27]
port 96 nsew signal tristate
flabel metal2 s 60032 79200 60144 80000 0 FreeSans 448 90 0 0 io_out[28]
port 97 nsew signal tristate
flabel metal2 s 62048 79200 62160 80000 0 FreeSans 448 90 0 0 io_out[29]
port 98 nsew signal tristate
flabel metal2 s 7616 79200 7728 80000 0 FreeSans 448 90 0 0 io_out[2]
port 99 nsew signal tristate
flabel metal2 s 64064 79200 64176 80000 0 FreeSans 448 90 0 0 io_out[30]
port 100 nsew signal tristate
flabel metal2 s 66080 79200 66192 80000 0 FreeSans 448 90 0 0 io_out[31]
port 101 nsew signal tristate
flabel metal2 s 68096 79200 68208 80000 0 FreeSans 448 90 0 0 io_out[32]
port 102 nsew signal tristate
flabel metal2 s 70112 79200 70224 80000 0 FreeSans 448 90 0 0 io_out[33]
port 103 nsew signal tristate
flabel metal2 s 72128 79200 72240 80000 0 FreeSans 448 90 0 0 io_out[34]
port 104 nsew signal tristate
flabel metal2 s 74144 79200 74256 80000 0 FreeSans 448 90 0 0 io_out[35]
port 105 nsew signal tristate
flabel metal2 s 76160 79200 76272 80000 0 FreeSans 448 90 0 0 io_out[36]
port 106 nsew signal tristate
flabel metal2 s 78176 79200 78288 80000 0 FreeSans 448 90 0 0 io_out[37]
port 107 nsew signal tristate
flabel metal2 s 9632 79200 9744 80000 0 FreeSans 448 90 0 0 io_out[3]
port 108 nsew signal tristate
flabel metal2 s 11648 79200 11760 80000 0 FreeSans 448 90 0 0 io_out[4]
port 109 nsew signal tristate
flabel metal2 s 13664 79200 13776 80000 0 FreeSans 448 90 0 0 io_out[5]
port 110 nsew signal tristate
flabel metal2 s 15680 79200 15792 80000 0 FreeSans 448 90 0 0 io_out[6]
port 111 nsew signal tristate
flabel metal2 s 17696 79200 17808 80000 0 FreeSans 448 90 0 0 io_out[7]
port 112 nsew signal tristate
flabel metal2 s 19712 79200 19824 80000 0 FreeSans 448 90 0 0 io_out[8]
port 113 nsew signal tristate
flabel metal2 s 21728 79200 21840 80000 0 FreeSans 448 90 0 0 io_out[9]
port 114 nsew signal tristate
flabel metal2 s 73024 0 73136 800 0 FreeSans 448 90 0 0 irq[0]
port 115 nsew signal tristate
flabel metal2 s 73248 0 73360 800 0 FreeSans 448 90 0 0 irq[1]
port 116 nsew signal tristate
flabel metal2 s 73472 0 73584 800 0 FreeSans 448 90 0 0 irq[2]
port 117 nsew signal tristate
flabel metal2 s 30016 0 30128 800 0 FreeSans 448 90 0 0 la_data_in[0]
port 118 nsew signal input
flabel metal2 s 36736 0 36848 800 0 FreeSans 448 90 0 0 la_data_in[10]
port 119 nsew signal input
flabel metal2 s 37408 0 37520 800 0 FreeSans 448 90 0 0 la_data_in[11]
port 120 nsew signal input
flabel metal2 s 38080 0 38192 800 0 FreeSans 448 90 0 0 la_data_in[12]
port 121 nsew signal input
flabel metal2 s 38752 0 38864 800 0 FreeSans 448 90 0 0 la_data_in[13]
port 122 nsew signal input
flabel metal2 s 39424 0 39536 800 0 FreeSans 448 90 0 0 la_data_in[14]
port 123 nsew signal input
flabel metal2 s 40096 0 40208 800 0 FreeSans 448 90 0 0 la_data_in[15]
port 124 nsew signal input
flabel metal2 s 40768 0 40880 800 0 FreeSans 448 90 0 0 la_data_in[16]
port 125 nsew signal input
flabel metal2 s 41440 0 41552 800 0 FreeSans 448 90 0 0 la_data_in[17]
port 126 nsew signal input
flabel metal2 s 42112 0 42224 800 0 FreeSans 448 90 0 0 la_data_in[18]
port 127 nsew signal input
flabel metal2 s 42784 0 42896 800 0 FreeSans 448 90 0 0 la_data_in[19]
port 128 nsew signal input
flabel metal2 s 30688 0 30800 800 0 FreeSans 448 90 0 0 la_data_in[1]
port 129 nsew signal input
flabel metal2 s 43456 0 43568 800 0 FreeSans 448 90 0 0 la_data_in[20]
port 130 nsew signal input
flabel metal2 s 44128 0 44240 800 0 FreeSans 448 90 0 0 la_data_in[21]
port 131 nsew signal input
flabel metal2 s 44800 0 44912 800 0 FreeSans 448 90 0 0 la_data_in[22]
port 132 nsew signal input
flabel metal2 s 45472 0 45584 800 0 FreeSans 448 90 0 0 la_data_in[23]
port 133 nsew signal input
flabel metal2 s 46144 0 46256 800 0 FreeSans 448 90 0 0 la_data_in[24]
port 134 nsew signal input
flabel metal2 s 46816 0 46928 800 0 FreeSans 448 90 0 0 la_data_in[25]
port 135 nsew signal input
flabel metal2 s 47488 0 47600 800 0 FreeSans 448 90 0 0 la_data_in[26]
port 136 nsew signal input
flabel metal2 s 48160 0 48272 800 0 FreeSans 448 90 0 0 la_data_in[27]
port 137 nsew signal input
flabel metal2 s 48832 0 48944 800 0 FreeSans 448 90 0 0 la_data_in[28]
port 138 nsew signal input
flabel metal2 s 49504 0 49616 800 0 FreeSans 448 90 0 0 la_data_in[29]
port 139 nsew signal input
flabel metal2 s 31360 0 31472 800 0 FreeSans 448 90 0 0 la_data_in[2]
port 140 nsew signal input
flabel metal2 s 50176 0 50288 800 0 FreeSans 448 90 0 0 la_data_in[30]
port 141 nsew signal input
flabel metal2 s 50848 0 50960 800 0 FreeSans 448 90 0 0 la_data_in[31]
port 142 nsew signal input
flabel metal2 s 51520 0 51632 800 0 FreeSans 448 90 0 0 la_data_in[32]
port 143 nsew signal input
flabel metal2 s 52192 0 52304 800 0 FreeSans 448 90 0 0 la_data_in[33]
port 144 nsew signal input
flabel metal2 s 52864 0 52976 800 0 FreeSans 448 90 0 0 la_data_in[34]
port 145 nsew signal input
flabel metal2 s 53536 0 53648 800 0 FreeSans 448 90 0 0 la_data_in[35]
port 146 nsew signal input
flabel metal2 s 54208 0 54320 800 0 FreeSans 448 90 0 0 la_data_in[36]
port 147 nsew signal input
flabel metal2 s 54880 0 54992 800 0 FreeSans 448 90 0 0 la_data_in[37]
port 148 nsew signal input
flabel metal2 s 55552 0 55664 800 0 FreeSans 448 90 0 0 la_data_in[38]
port 149 nsew signal input
flabel metal2 s 56224 0 56336 800 0 FreeSans 448 90 0 0 la_data_in[39]
port 150 nsew signal input
flabel metal2 s 32032 0 32144 800 0 FreeSans 448 90 0 0 la_data_in[3]
port 151 nsew signal input
flabel metal2 s 56896 0 57008 800 0 FreeSans 448 90 0 0 la_data_in[40]
port 152 nsew signal input
flabel metal2 s 57568 0 57680 800 0 FreeSans 448 90 0 0 la_data_in[41]
port 153 nsew signal input
flabel metal2 s 58240 0 58352 800 0 FreeSans 448 90 0 0 la_data_in[42]
port 154 nsew signal input
flabel metal2 s 58912 0 59024 800 0 FreeSans 448 90 0 0 la_data_in[43]
port 155 nsew signal input
flabel metal2 s 59584 0 59696 800 0 FreeSans 448 90 0 0 la_data_in[44]
port 156 nsew signal input
flabel metal2 s 60256 0 60368 800 0 FreeSans 448 90 0 0 la_data_in[45]
port 157 nsew signal input
flabel metal2 s 60928 0 61040 800 0 FreeSans 448 90 0 0 la_data_in[46]
port 158 nsew signal input
flabel metal2 s 61600 0 61712 800 0 FreeSans 448 90 0 0 la_data_in[47]
port 159 nsew signal input
flabel metal2 s 62272 0 62384 800 0 FreeSans 448 90 0 0 la_data_in[48]
port 160 nsew signal input
flabel metal2 s 62944 0 63056 800 0 FreeSans 448 90 0 0 la_data_in[49]
port 161 nsew signal input
flabel metal2 s 32704 0 32816 800 0 FreeSans 448 90 0 0 la_data_in[4]
port 162 nsew signal input
flabel metal2 s 63616 0 63728 800 0 FreeSans 448 90 0 0 la_data_in[50]
port 163 nsew signal input
flabel metal2 s 64288 0 64400 800 0 FreeSans 448 90 0 0 la_data_in[51]
port 164 nsew signal input
flabel metal2 s 64960 0 65072 800 0 FreeSans 448 90 0 0 la_data_in[52]
port 165 nsew signal input
flabel metal2 s 65632 0 65744 800 0 FreeSans 448 90 0 0 la_data_in[53]
port 166 nsew signal input
flabel metal2 s 66304 0 66416 800 0 FreeSans 448 90 0 0 la_data_in[54]
port 167 nsew signal input
flabel metal2 s 66976 0 67088 800 0 FreeSans 448 90 0 0 la_data_in[55]
port 168 nsew signal input
flabel metal2 s 67648 0 67760 800 0 FreeSans 448 90 0 0 la_data_in[56]
port 169 nsew signal input
flabel metal2 s 68320 0 68432 800 0 FreeSans 448 90 0 0 la_data_in[57]
port 170 nsew signal input
flabel metal2 s 68992 0 69104 800 0 FreeSans 448 90 0 0 la_data_in[58]
port 171 nsew signal input
flabel metal2 s 69664 0 69776 800 0 FreeSans 448 90 0 0 la_data_in[59]
port 172 nsew signal input
flabel metal2 s 33376 0 33488 800 0 FreeSans 448 90 0 0 la_data_in[5]
port 173 nsew signal input
flabel metal2 s 70336 0 70448 800 0 FreeSans 448 90 0 0 la_data_in[60]
port 174 nsew signal input
flabel metal2 s 71008 0 71120 800 0 FreeSans 448 90 0 0 la_data_in[61]
port 175 nsew signal input
flabel metal2 s 71680 0 71792 800 0 FreeSans 448 90 0 0 la_data_in[62]
port 176 nsew signal input
flabel metal2 s 72352 0 72464 800 0 FreeSans 448 90 0 0 la_data_in[63]
port 177 nsew signal input
flabel metal2 s 34048 0 34160 800 0 FreeSans 448 90 0 0 la_data_in[6]
port 178 nsew signal input
flabel metal2 s 34720 0 34832 800 0 FreeSans 448 90 0 0 la_data_in[7]
port 179 nsew signal input
flabel metal2 s 35392 0 35504 800 0 FreeSans 448 90 0 0 la_data_in[8]
port 180 nsew signal input
flabel metal2 s 36064 0 36176 800 0 FreeSans 448 90 0 0 la_data_in[9]
port 181 nsew signal input
flabel metal2 s 30240 0 30352 800 0 FreeSans 448 90 0 0 la_data_out[0]
port 182 nsew signal tristate
flabel metal2 s 36960 0 37072 800 0 FreeSans 448 90 0 0 la_data_out[10]
port 183 nsew signal tristate
flabel metal2 s 37632 0 37744 800 0 FreeSans 448 90 0 0 la_data_out[11]
port 184 nsew signal tristate
flabel metal2 s 38304 0 38416 800 0 FreeSans 448 90 0 0 la_data_out[12]
port 185 nsew signal tristate
flabel metal2 s 38976 0 39088 800 0 FreeSans 448 90 0 0 la_data_out[13]
port 186 nsew signal tristate
flabel metal2 s 39648 0 39760 800 0 FreeSans 448 90 0 0 la_data_out[14]
port 187 nsew signal tristate
flabel metal2 s 40320 0 40432 800 0 FreeSans 448 90 0 0 la_data_out[15]
port 188 nsew signal tristate
flabel metal2 s 40992 0 41104 800 0 FreeSans 448 90 0 0 la_data_out[16]
port 189 nsew signal tristate
flabel metal2 s 41664 0 41776 800 0 FreeSans 448 90 0 0 la_data_out[17]
port 190 nsew signal tristate
flabel metal2 s 42336 0 42448 800 0 FreeSans 448 90 0 0 la_data_out[18]
port 191 nsew signal tristate
flabel metal2 s 43008 0 43120 800 0 FreeSans 448 90 0 0 la_data_out[19]
port 192 nsew signal tristate
flabel metal2 s 30912 0 31024 800 0 FreeSans 448 90 0 0 la_data_out[1]
port 193 nsew signal tristate
flabel metal2 s 43680 0 43792 800 0 FreeSans 448 90 0 0 la_data_out[20]
port 194 nsew signal tristate
flabel metal2 s 44352 0 44464 800 0 FreeSans 448 90 0 0 la_data_out[21]
port 195 nsew signal tristate
flabel metal2 s 45024 0 45136 800 0 FreeSans 448 90 0 0 la_data_out[22]
port 196 nsew signal tristate
flabel metal2 s 45696 0 45808 800 0 FreeSans 448 90 0 0 la_data_out[23]
port 197 nsew signal tristate
flabel metal2 s 46368 0 46480 800 0 FreeSans 448 90 0 0 la_data_out[24]
port 198 nsew signal tristate
flabel metal2 s 47040 0 47152 800 0 FreeSans 448 90 0 0 la_data_out[25]
port 199 nsew signal tristate
flabel metal2 s 47712 0 47824 800 0 FreeSans 448 90 0 0 la_data_out[26]
port 200 nsew signal tristate
flabel metal2 s 48384 0 48496 800 0 FreeSans 448 90 0 0 la_data_out[27]
port 201 nsew signal tristate
flabel metal2 s 49056 0 49168 800 0 FreeSans 448 90 0 0 la_data_out[28]
port 202 nsew signal tristate
flabel metal2 s 49728 0 49840 800 0 FreeSans 448 90 0 0 la_data_out[29]
port 203 nsew signal tristate
flabel metal2 s 31584 0 31696 800 0 FreeSans 448 90 0 0 la_data_out[2]
port 204 nsew signal tristate
flabel metal2 s 50400 0 50512 800 0 FreeSans 448 90 0 0 la_data_out[30]
port 205 nsew signal tristate
flabel metal2 s 51072 0 51184 800 0 FreeSans 448 90 0 0 la_data_out[31]
port 206 nsew signal tristate
flabel metal2 s 51744 0 51856 800 0 FreeSans 448 90 0 0 la_data_out[32]
port 207 nsew signal tristate
flabel metal2 s 52416 0 52528 800 0 FreeSans 448 90 0 0 la_data_out[33]
port 208 nsew signal tristate
flabel metal2 s 53088 0 53200 800 0 FreeSans 448 90 0 0 la_data_out[34]
port 209 nsew signal tristate
flabel metal2 s 53760 0 53872 800 0 FreeSans 448 90 0 0 la_data_out[35]
port 210 nsew signal tristate
flabel metal2 s 54432 0 54544 800 0 FreeSans 448 90 0 0 la_data_out[36]
port 211 nsew signal tristate
flabel metal2 s 55104 0 55216 800 0 FreeSans 448 90 0 0 la_data_out[37]
port 212 nsew signal tristate
flabel metal2 s 55776 0 55888 800 0 FreeSans 448 90 0 0 la_data_out[38]
port 213 nsew signal tristate
flabel metal2 s 56448 0 56560 800 0 FreeSans 448 90 0 0 la_data_out[39]
port 214 nsew signal tristate
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 la_data_out[3]
port 215 nsew signal tristate
flabel metal2 s 57120 0 57232 800 0 FreeSans 448 90 0 0 la_data_out[40]
port 216 nsew signal tristate
flabel metal2 s 57792 0 57904 800 0 FreeSans 448 90 0 0 la_data_out[41]
port 217 nsew signal tristate
flabel metal2 s 58464 0 58576 800 0 FreeSans 448 90 0 0 la_data_out[42]
port 218 nsew signal tristate
flabel metal2 s 59136 0 59248 800 0 FreeSans 448 90 0 0 la_data_out[43]
port 219 nsew signal tristate
flabel metal2 s 59808 0 59920 800 0 FreeSans 448 90 0 0 la_data_out[44]
port 220 nsew signal tristate
flabel metal2 s 60480 0 60592 800 0 FreeSans 448 90 0 0 la_data_out[45]
port 221 nsew signal tristate
flabel metal2 s 61152 0 61264 800 0 FreeSans 448 90 0 0 la_data_out[46]
port 222 nsew signal tristate
flabel metal2 s 61824 0 61936 800 0 FreeSans 448 90 0 0 la_data_out[47]
port 223 nsew signal tristate
flabel metal2 s 62496 0 62608 800 0 FreeSans 448 90 0 0 la_data_out[48]
port 224 nsew signal tristate
flabel metal2 s 63168 0 63280 800 0 FreeSans 448 90 0 0 la_data_out[49]
port 225 nsew signal tristate
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 la_data_out[4]
port 226 nsew signal tristate
flabel metal2 s 63840 0 63952 800 0 FreeSans 448 90 0 0 la_data_out[50]
port 227 nsew signal tristate
flabel metal2 s 64512 0 64624 800 0 FreeSans 448 90 0 0 la_data_out[51]
port 228 nsew signal tristate
flabel metal2 s 65184 0 65296 800 0 FreeSans 448 90 0 0 la_data_out[52]
port 229 nsew signal tristate
flabel metal2 s 65856 0 65968 800 0 FreeSans 448 90 0 0 la_data_out[53]
port 230 nsew signal tristate
flabel metal2 s 66528 0 66640 800 0 FreeSans 448 90 0 0 la_data_out[54]
port 231 nsew signal tristate
flabel metal2 s 67200 0 67312 800 0 FreeSans 448 90 0 0 la_data_out[55]
port 232 nsew signal tristate
flabel metal2 s 67872 0 67984 800 0 FreeSans 448 90 0 0 la_data_out[56]
port 233 nsew signal tristate
flabel metal2 s 68544 0 68656 800 0 FreeSans 448 90 0 0 la_data_out[57]
port 234 nsew signal tristate
flabel metal2 s 69216 0 69328 800 0 FreeSans 448 90 0 0 la_data_out[58]
port 235 nsew signal tristate
flabel metal2 s 69888 0 70000 800 0 FreeSans 448 90 0 0 la_data_out[59]
port 236 nsew signal tristate
flabel metal2 s 33600 0 33712 800 0 FreeSans 448 90 0 0 la_data_out[5]
port 237 nsew signal tristate
flabel metal2 s 70560 0 70672 800 0 FreeSans 448 90 0 0 la_data_out[60]
port 238 nsew signal tristate
flabel metal2 s 71232 0 71344 800 0 FreeSans 448 90 0 0 la_data_out[61]
port 239 nsew signal tristate
flabel metal2 s 71904 0 72016 800 0 FreeSans 448 90 0 0 la_data_out[62]
port 240 nsew signal tristate
flabel metal2 s 72576 0 72688 800 0 FreeSans 448 90 0 0 la_data_out[63]
port 241 nsew signal tristate
flabel metal2 s 34272 0 34384 800 0 FreeSans 448 90 0 0 la_data_out[6]
port 242 nsew signal tristate
flabel metal2 s 34944 0 35056 800 0 FreeSans 448 90 0 0 la_data_out[7]
port 243 nsew signal tristate
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 la_data_out[8]
port 244 nsew signal tristate
flabel metal2 s 36288 0 36400 800 0 FreeSans 448 90 0 0 la_data_out[9]
port 245 nsew signal tristate
flabel metal2 s 30464 0 30576 800 0 FreeSans 448 90 0 0 la_oenb[0]
port 246 nsew signal input
flabel metal2 s 37184 0 37296 800 0 FreeSans 448 90 0 0 la_oenb[10]
port 247 nsew signal input
flabel metal2 s 37856 0 37968 800 0 FreeSans 448 90 0 0 la_oenb[11]
port 248 nsew signal input
flabel metal2 s 38528 0 38640 800 0 FreeSans 448 90 0 0 la_oenb[12]
port 249 nsew signal input
flabel metal2 s 39200 0 39312 800 0 FreeSans 448 90 0 0 la_oenb[13]
port 250 nsew signal input
flabel metal2 s 39872 0 39984 800 0 FreeSans 448 90 0 0 la_oenb[14]
port 251 nsew signal input
flabel metal2 s 40544 0 40656 800 0 FreeSans 448 90 0 0 la_oenb[15]
port 252 nsew signal input
flabel metal2 s 41216 0 41328 800 0 FreeSans 448 90 0 0 la_oenb[16]
port 253 nsew signal input
flabel metal2 s 41888 0 42000 800 0 FreeSans 448 90 0 0 la_oenb[17]
port 254 nsew signal input
flabel metal2 s 42560 0 42672 800 0 FreeSans 448 90 0 0 la_oenb[18]
port 255 nsew signal input
flabel metal2 s 43232 0 43344 800 0 FreeSans 448 90 0 0 la_oenb[19]
port 256 nsew signal input
flabel metal2 s 31136 0 31248 800 0 FreeSans 448 90 0 0 la_oenb[1]
port 257 nsew signal input
flabel metal2 s 43904 0 44016 800 0 FreeSans 448 90 0 0 la_oenb[20]
port 258 nsew signal input
flabel metal2 s 44576 0 44688 800 0 FreeSans 448 90 0 0 la_oenb[21]
port 259 nsew signal input
flabel metal2 s 45248 0 45360 800 0 FreeSans 448 90 0 0 la_oenb[22]
port 260 nsew signal input
flabel metal2 s 45920 0 46032 800 0 FreeSans 448 90 0 0 la_oenb[23]
port 261 nsew signal input
flabel metal2 s 46592 0 46704 800 0 FreeSans 448 90 0 0 la_oenb[24]
port 262 nsew signal input
flabel metal2 s 47264 0 47376 800 0 FreeSans 448 90 0 0 la_oenb[25]
port 263 nsew signal input
flabel metal2 s 47936 0 48048 800 0 FreeSans 448 90 0 0 la_oenb[26]
port 264 nsew signal input
flabel metal2 s 48608 0 48720 800 0 FreeSans 448 90 0 0 la_oenb[27]
port 265 nsew signal input
flabel metal2 s 49280 0 49392 800 0 FreeSans 448 90 0 0 la_oenb[28]
port 266 nsew signal input
flabel metal2 s 49952 0 50064 800 0 FreeSans 448 90 0 0 la_oenb[29]
port 267 nsew signal input
flabel metal2 s 31808 0 31920 800 0 FreeSans 448 90 0 0 la_oenb[2]
port 268 nsew signal input
flabel metal2 s 50624 0 50736 800 0 FreeSans 448 90 0 0 la_oenb[30]
port 269 nsew signal input
flabel metal2 s 51296 0 51408 800 0 FreeSans 448 90 0 0 la_oenb[31]
port 270 nsew signal input
flabel metal2 s 51968 0 52080 800 0 FreeSans 448 90 0 0 la_oenb[32]
port 271 nsew signal input
flabel metal2 s 52640 0 52752 800 0 FreeSans 448 90 0 0 la_oenb[33]
port 272 nsew signal input
flabel metal2 s 53312 0 53424 800 0 FreeSans 448 90 0 0 la_oenb[34]
port 273 nsew signal input
flabel metal2 s 53984 0 54096 800 0 FreeSans 448 90 0 0 la_oenb[35]
port 274 nsew signal input
flabel metal2 s 54656 0 54768 800 0 FreeSans 448 90 0 0 la_oenb[36]
port 275 nsew signal input
flabel metal2 s 55328 0 55440 800 0 FreeSans 448 90 0 0 la_oenb[37]
port 276 nsew signal input
flabel metal2 s 56000 0 56112 800 0 FreeSans 448 90 0 0 la_oenb[38]
port 277 nsew signal input
flabel metal2 s 56672 0 56784 800 0 FreeSans 448 90 0 0 la_oenb[39]
port 278 nsew signal input
flabel metal2 s 32480 0 32592 800 0 FreeSans 448 90 0 0 la_oenb[3]
port 279 nsew signal input
flabel metal2 s 57344 0 57456 800 0 FreeSans 448 90 0 0 la_oenb[40]
port 280 nsew signal input
flabel metal2 s 58016 0 58128 800 0 FreeSans 448 90 0 0 la_oenb[41]
port 281 nsew signal input
flabel metal2 s 58688 0 58800 800 0 FreeSans 448 90 0 0 la_oenb[42]
port 282 nsew signal input
flabel metal2 s 59360 0 59472 800 0 FreeSans 448 90 0 0 la_oenb[43]
port 283 nsew signal input
flabel metal2 s 60032 0 60144 800 0 FreeSans 448 90 0 0 la_oenb[44]
port 284 nsew signal input
flabel metal2 s 60704 0 60816 800 0 FreeSans 448 90 0 0 la_oenb[45]
port 285 nsew signal input
flabel metal2 s 61376 0 61488 800 0 FreeSans 448 90 0 0 la_oenb[46]
port 286 nsew signal input
flabel metal2 s 62048 0 62160 800 0 FreeSans 448 90 0 0 la_oenb[47]
port 287 nsew signal input
flabel metal2 s 62720 0 62832 800 0 FreeSans 448 90 0 0 la_oenb[48]
port 288 nsew signal input
flabel metal2 s 63392 0 63504 800 0 FreeSans 448 90 0 0 la_oenb[49]
port 289 nsew signal input
flabel metal2 s 33152 0 33264 800 0 FreeSans 448 90 0 0 la_oenb[4]
port 290 nsew signal input
flabel metal2 s 64064 0 64176 800 0 FreeSans 448 90 0 0 la_oenb[50]
port 291 nsew signal input
flabel metal2 s 64736 0 64848 800 0 FreeSans 448 90 0 0 la_oenb[51]
port 292 nsew signal input
flabel metal2 s 65408 0 65520 800 0 FreeSans 448 90 0 0 la_oenb[52]
port 293 nsew signal input
flabel metal2 s 66080 0 66192 800 0 FreeSans 448 90 0 0 la_oenb[53]
port 294 nsew signal input
flabel metal2 s 66752 0 66864 800 0 FreeSans 448 90 0 0 la_oenb[54]
port 295 nsew signal input
flabel metal2 s 67424 0 67536 800 0 FreeSans 448 90 0 0 la_oenb[55]
port 296 nsew signal input
flabel metal2 s 68096 0 68208 800 0 FreeSans 448 90 0 0 la_oenb[56]
port 297 nsew signal input
flabel metal2 s 68768 0 68880 800 0 FreeSans 448 90 0 0 la_oenb[57]
port 298 nsew signal input
flabel metal2 s 69440 0 69552 800 0 FreeSans 448 90 0 0 la_oenb[58]
port 299 nsew signal input
flabel metal2 s 70112 0 70224 800 0 FreeSans 448 90 0 0 la_oenb[59]
port 300 nsew signal input
flabel metal2 s 33824 0 33936 800 0 FreeSans 448 90 0 0 la_oenb[5]
port 301 nsew signal input
flabel metal2 s 70784 0 70896 800 0 FreeSans 448 90 0 0 la_oenb[60]
port 302 nsew signal input
flabel metal2 s 71456 0 71568 800 0 FreeSans 448 90 0 0 la_oenb[61]
port 303 nsew signal input
flabel metal2 s 72128 0 72240 800 0 FreeSans 448 90 0 0 la_oenb[62]
port 304 nsew signal input
flabel metal2 s 72800 0 72912 800 0 FreeSans 448 90 0 0 la_oenb[63]
port 305 nsew signal input
flabel metal2 s 34496 0 34608 800 0 FreeSans 448 90 0 0 la_oenb[6]
port 306 nsew signal input
flabel metal2 s 35168 0 35280 800 0 FreeSans 448 90 0 0 la_oenb[7]
port 307 nsew signal input
flabel metal2 s 35840 0 35952 800 0 FreeSans 448 90 0 0 la_oenb[8]
port 308 nsew signal input
flabel metal2 s 36512 0 36624 800 0 FreeSans 448 90 0 0 la_oenb[9]
port 309 nsew signal input
flabel metal4 s 4448 3076 4768 76892 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 35168 3076 35488 76892 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 65888 3076 66208 76892 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 19808 3076 20128 76892 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 76892 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 6272 0 6384 800 0 FreeSans 448 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 6496 0 6608 800 0 FreeSans 448 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 7616 0 7728 800 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 15232 0 15344 800 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 15904 0 16016 800 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 16576 0 16688 800 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 17248 0 17360 800 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 17920 0 18032 800 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 18592 0 18704 800 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 19264 0 19376 800 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 19936 0 20048 800 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 20608 0 20720 800 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 21280 0 21392 800 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 8512 0 8624 800 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 21952 0 22064 800 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 22624 0 22736 800 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 23296 0 23408 800 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 23968 0 24080 800 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 24640 0 24752 800 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 25312 0 25424 800 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 25984 0 26096 800 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 26656 0 26768 800 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 27328 0 27440 800 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 28000 0 28112 800 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 28672 0 28784 800 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 29344 0 29456 800 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 10304 0 10416 800 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 11200 0 11312 800 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 11872 0 11984 800 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 12544 0 12656 800 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 13216 0 13328 800 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 13888 0 14000 800 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 14560 0 14672 800 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 6944 0 7056 800 0 FreeSans 448 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 7840 0 7952 800 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 27552 0 27664 800 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 28224 0 28336 800 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 9632 0 9744 800 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 10528 0 10640 800 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 11424 0 11536 800 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 12768 0 12880 800 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 14112 0 14224 800 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 15680 0 15792 800 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 16352 0 16464 800 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 17024 0 17136 800 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 17696 0 17808 800 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 18368 0 18480 800 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 19040 0 19152 800 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 19712 0 19824 800 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 20384 0 20496 800 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 21056 0 21168 800 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 21728 0 21840 800 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 8960 0 9072 800 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 22400 0 22512 800 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 23072 0 23184 800 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 23744 0 23856 800 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 24416 0 24528 800 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 25088 0 25200 800 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 25760 0 25872 800 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 26432 0 26544 800 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 27104 0 27216 800 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 27776 0 27888 800 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 28448 0 28560 800 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 9856 0 9968 800 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 29120 0 29232 800 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 29792 0 29904 800 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 11648 0 11760 800 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 12320 0 12432 800 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 12992 0 13104 800 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 13664 0 13776 800 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 14336 0 14448 800 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 15008 0 15120 800 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 8288 0 8400 800 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 9184 0 9296 800 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 10976 0 11088 800 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 7168 0 7280 800 0 FreeSans 448 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel metal1 39984 76048 39984 76048 0 vdd
rlabel metal1 39984 76832 39984 76832 0 vss
rlabel metal2 39480 75656 39480 75656 0 _000_
rlabel metal2 41664 75096 41664 75096 0 _001_
rlabel metal2 37800 72744 37800 72744 0 _002_
rlabel metal2 39816 75376 39816 75376 0 _003_
rlabel metal2 31192 75096 31192 75096 0 _004_
rlabel metal2 53704 75600 53704 75600 0 _005_
rlabel metal3 55552 75768 55552 75768 0 _006_
rlabel metal2 56056 72912 56056 72912 0 _007_
rlabel metal2 55384 75152 55384 75152 0 _008_
rlabel metal2 30184 75544 30184 75544 0 _009_
rlabel metal2 30464 75656 30464 75656 0 _010_
rlabel metal2 29344 75544 29344 75544 0 _011_
rlabel metal2 30072 75264 30072 75264 0 _012_
rlabel metal2 31416 73584 31416 73584 0 _013_
rlabel metal3 37912 73304 37912 73304 0 _014_
rlabel metal2 36680 72464 36680 72464 0 _015_
rlabel metal3 37016 72408 37016 72408 0 _016_
rlabel metal2 36736 72744 36736 72744 0 _017_
rlabel metal2 40432 73528 40432 73528 0 _018_
rlabel metal2 34104 75152 34104 75152 0 _019_
rlabel metal2 58688 71848 58688 71848 0 _020_
rlabel metal3 58352 73528 58352 73528 0 _021_
rlabel metal3 59472 73976 59472 73976 0 _022_
rlabel metal2 60312 74368 60312 74368 0 _023_
rlabel metal3 52696 75488 52696 75488 0 _024_
rlabel metal2 34440 76608 34440 76608 0 _025_
rlabel metal2 33880 73584 33880 73584 0 _026_
rlabel metal2 32256 75096 32256 75096 0 _027_
rlabel metal3 33040 74200 33040 74200 0 _028_
rlabel metal2 41944 70952 41944 70952 0 _029_
rlabel metal2 40600 74536 40600 74536 0 _030_
rlabel metal2 42840 74480 42840 74480 0 _031_
rlabel metal3 43512 74088 43512 74088 0 _032_
rlabel metal2 35616 74088 35616 74088 0 _033_
rlabel metal2 52696 73304 52696 73304 0 _034_
rlabel metal2 51072 75656 51072 75656 0 _035_
rlabel metal2 54264 74648 54264 74648 0 _036_
rlabel metal2 54488 73752 54488 73752 0 _037_
rlabel metal2 54264 76440 54264 76440 0 _038_
rlabel metal3 36792 74088 36792 74088 0 _039_
rlabel metal3 35056 73976 35056 73976 0 _040_
rlabel metal2 42784 70392 42784 70392 0 _041_
rlabel metal2 38360 72912 38360 72912 0 _042_
rlabel metal3 38640 73528 38640 73528 0 _043_
rlabel metal2 36568 74200 36568 74200 0 _044_
rlabel metal2 36904 74368 36904 74368 0 _045_
rlabel metal2 36456 75096 36456 75096 0 _046_
rlabel metal3 51464 71736 51464 71736 0 _047_
rlabel metal2 49952 73416 49952 73416 0 _048_
rlabel metal3 49448 76552 49448 76552 0 _049_
rlabel metal2 49672 76104 49672 76104 0 _050_
rlabel metal2 47880 75544 47880 75544 0 _051_
rlabel metal2 36120 75824 36120 75824 0 _052_
rlabel metal2 50008 75656 50008 75656 0 _053_
rlabel metal2 30408 72968 30408 72968 0 _054_
rlabel metal2 38024 73864 38024 73864 0 _055_
rlabel metal2 38024 74368 38024 74368 0 _056_
rlabel metal2 29400 74592 29400 74592 0 _057_
rlabel metal2 35336 75320 35336 75320 0 _058_
rlabel metal2 46872 75096 46872 75096 0 _059_
rlabel metal2 43288 75040 43288 75040 0 _060_
rlabel metal2 42224 75432 42224 75432 0 _061_
rlabel metal2 46312 70504 46312 70504 0 _062_
rlabel metal3 45976 73416 45976 73416 0 _063_
rlabel metal2 45640 72632 45640 72632 0 _064_
rlabel metal2 44184 72072 44184 72072 0 _065_
rlabel metal2 42616 72856 42616 72856 0 _066_
rlabel metal3 46536 73528 46536 73528 0 _067_
rlabel metal2 46312 73528 46312 73528 0 _068_
rlabel metal2 43960 70504 43960 70504 0 _069_
rlabel metal2 43008 71736 43008 71736 0 _070_
rlabel metal2 39144 72128 39144 72128 0 _071_
rlabel metal2 37688 72240 37688 72240 0 _072_
rlabel metal2 45752 72632 45752 72632 0 _073_
rlabel metal3 39256 71176 39256 71176 0 _074_
rlabel metal2 39200 71176 39200 71176 0 _075_
rlabel metal3 38752 70168 38752 70168 0 _076_
rlabel metal2 38696 73472 38696 73472 0 _077_
rlabel metal2 40264 72520 40264 72520 0 _078_
rlabel metal3 40656 71064 40656 71064 0 _079_
rlabel metal2 43568 70392 43568 70392 0 _080_
rlabel metal2 43848 72128 43848 72128 0 _081_
rlabel metal2 45528 71736 45528 71736 0 _082_
rlabel metal3 44744 72520 44744 72520 0 _083_
rlabel metal2 43568 73304 43568 73304 0 _084_
rlabel metal2 44072 73864 44072 73864 0 _085_
rlabel metal2 43512 76160 43512 76160 0 _086_
rlabel metal3 58744 74984 58744 74984 0 _087_
rlabel metal2 54376 74928 54376 74928 0 _088_
rlabel metal3 54208 73976 54208 73976 0 _089_
rlabel metal3 52360 73864 52360 73864 0 _090_
rlabel metal3 56616 75432 56616 75432 0 _091_
rlabel metal3 52024 75432 52024 75432 0 _092_
rlabel metal2 52192 74088 52192 74088 0 _093_
rlabel metal2 51800 72520 51800 72520 0 _094_
rlabel metal3 49168 73192 49168 73192 0 _095_
rlabel metal2 59640 73416 59640 73416 0 _096_
rlabel metal2 59304 73528 59304 73528 0 _097_
rlabel metal2 54320 71736 54320 71736 0 _098_
rlabel metal3 52360 72520 52360 72520 0 _099_
rlabel metal3 58184 72520 58184 72520 0 _100_
rlabel metal2 57624 73696 57624 73696 0 _101_
rlabel metal3 58688 73416 58688 73416 0 _102_
rlabel metal2 57512 72800 57512 72800 0 _103_
rlabel metal2 56616 72296 56616 72296 0 _104_
rlabel metal2 57288 74088 57288 74088 0 _105_
rlabel metal2 58072 72632 58072 72632 0 _106_
rlabel metal2 57848 72072 57848 72072 0 _107_
rlabel metal2 52472 72968 52472 72968 0 _108_
rlabel metal2 52920 72576 52920 72576 0 _109_
rlabel metal2 49896 73024 49896 73024 0 _110_
rlabel metal2 51184 73416 51184 73416 0 _111_
rlabel metal3 50568 73080 50568 73080 0 _112_
rlabel metal2 50512 73528 50512 73528 0 _113_
rlabel metal2 50120 72296 50120 72296 0 _114_
rlabel metal2 49840 74312 49840 74312 0 _115_
rlabel metal3 51184 73864 51184 73864 0 _116_
rlabel metal2 52584 75936 52584 75936 0 _117_
rlabel metal2 44968 71064 44968 71064 0 _118_
rlabel metal2 1792 76552 1792 76552 0 io_active
rlabel metal2 38584 75264 38584 75264 0 io_in[18]
rlabel metal2 40880 69496 40880 69496 0 io_in[19]
rlabel metal2 45528 70448 45528 70448 0 io_in[20]
rlabel metal3 45920 69496 45920 69496 0 io_in[21]
rlabel metal2 48328 71456 48328 71456 0 io_in[22]
rlabel metal2 48272 70392 48272 70392 0 io_in[23]
rlabel metal2 54824 76832 54824 76832 0 io_in[24]
rlabel metal2 52080 76440 52080 76440 0 io_in[25]
rlabel metal2 55048 75600 55048 75600 0 io_in[26]
rlabel metal3 57344 76552 57344 76552 0 io_in[27]
rlabel metal3 59024 76552 59024 76552 0 io_in[28]
rlabel metal2 61320 76832 61320 76832 0 io_in[29]
rlabel metal2 62832 73528 62832 73528 0 io_in[30]
rlabel metal2 65408 75096 65408 75096 0 io_in[31]
rlabel metal3 69664 75768 69664 75768 0 io_in[32]
rlabel metal3 69272 75432 69272 75432 0 io_in[33]
rlabel metal2 70840 77154 70840 77154 0 io_in[34]
rlabel metal2 73080 76440 73080 76440 0 io_in[35]
rlabel metal3 75488 75544 75488 75544 0 io_in[36]
rlabel metal3 77280 74984 77280 74984 0 io_in[37]
rlabel metal3 4760 76552 4760 76552 0 io_out[0]
rlabel metal2 23800 77770 23800 77770 0 io_out[10]
rlabel metal2 25816 77770 25816 77770 0 io_out[11]
rlabel metal2 27832 77770 27832 77770 0 io_out[12]
rlabel metal2 30184 77168 30184 77168 0 io_out[13]
rlabel metal2 31864 77490 31864 77490 0 io_out[14]
rlabel metal2 33936 76328 33936 76328 0 io_out[15]
rlabel metal2 35896 77770 35896 77770 0 io_out[16]
rlabel metal2 37912 78106 37912 78106 0 io_out[17]
rlabel metal2 11704 77882 11704 77882 0 io_out[4]
rlabel metal2 13776 76552 13776 76552 0 io_out[5]
rlabel metal2 15736 77770 15736 77770 0 io_out[6]
rlabel metal2 17752 77882 17752 77882 0 io_out[7]
rlabel metal2 19656 77056 19656 77056 0 io_out[8]
rlabel metal2 21840 76328 21840 76328 0 io_out[9]
rlabel metal2 3360 76328 3360 76328 0 net1
rlabel metal3 59472 75880 59472 75880 0 net10
rlabel metal2 7112 75544 7112 75544 0 net100
rlabel metal2 8960 76664 8960 76664 0 net101
rlabel metal2 11032 77938 11032 77938 0 net102
rlabel metal3 13384 75544 13384 75544 0 net103
rlabel metal2 15176 75544 15176 75544 0 net104
rlabel metal2 17192 75544 17192 75544 0 net105
rlabel metal2 19208 75544 19208 75544 0 net106
rlabel metal3 21392 75544 21392 75544 0 net107
rlabel metal2 23240 75544 23240 75544 0 net108
rlabel metal2 25256 75544 25256 75544 0 net109
rlabel metal2 56728 73136 56728 73136 0 net11
rlabel metal2 27160 77378 27160 77378 0 net110
rlabel metal3 28560 75544 28560 75544 0 net111
rlabel metal2 31640 74984 31640 74984 0 net112
rlabel metal2 29960 76048 29960 76048 0 net113
rlabel metal2 35448 72352 35448 72352 0 net114
rlabel metal2 36064 72408 36064 72408 0 net115
rlabel metal2 39032 72016 39032 72016 0 net116
rlabel metal2 41608 70560 41608 70560 0 net117
rlabel metal2 47768 73752 47768 73752 0 net118
rlabel metal3 47152 75432 47152 75432 0 net119
rlabel metal2 53928 73696 53928 73696 0 net12
rlabel metal2 47768 72856 47768 72856 0 net120
rlabel metal2 55832 76832 55832 76832 0 net121
rlabel metal2 51520 70840 51520 70840 0 net122
rlabel metal2 53648 70840 53648 70840 0 net123
rlabel metal2 55384 77938 55384 77938 0 net124
rlabel metal2 63224 76720 63224 76720 0 net125
rlabel metal3 60592 73864 60592 73864 0 net126
rlabel metal3 62048 75096 62048 75096 0 net127
rlabel metal3 63728 75096 63728 75096 0 net128
rlabel metal3 66080 75544 66080 75544 0 net129
rlabel metal2 54152 70616 54152 70616 0 net13
rlabel metal3 67760 75544 67760 75544 0 net130
rlabel metal3 69888 75544 69888 75544 0 net131
rlabel metal2 72408 76720 72408 76720 0 net132
rlabel metal3 74088 76664 74088 76664 0 net133
rlabel metal3 75936 76664 75936 76664 0 net134
rlabel metal2 77672 76664 77672 76664 0 net135
rlabel metal2 5768 75544 5768 75544 0 net136
rlabel metal2 7784 76664 7784 76664 0 net137
rlabel metal2 9800 76664 9800 76664 0 net138
rlabel metal2 35784 74312 35784 74312 0 net139
rlabel metal2 59976 75656 59976 75656 0 net14
rlabel metal2 47096 73808 47096 73808 0 net140
rlabel metal3 45752 74648 45752 74648 0 net141
rlabel metal2 46648 72352 46648 72352 0 net142
rlabel metal2 48384 72408 48384 72408 0 net143
rlabel metal2 49672 76776 49672 76776 0 net144
rlabel metal2 52248 72352 52248 72352 0 net145
rlabel metal2 54040 77378 54040 77378 0 net146
rlabel metal2 62552 76832 62552 76832 0 net147
rlabel metal2 61992 75152 61992 75152 0 net148
rlabel metal2 60872 73640 60872 73640 0 net149
rlabel metal2 55384 71568 55384 71568 0 net15
rlabel metal2 63336 75320 63336 75320 0 net150
rlabel metal3 65072 75432 65072 75432 0 net151
rlabel metal2 66360 75824 66360 75824 0 net152
rlabel metal2 68376 75264 68376 75264 0 net153
rlabel metal3 70840 76552 70840 76552 0 net154
rlabel metal2 73976 76776 73976 76776 0 net155
rlabel metal2 75320 76944 75320 76944 0 net156
rlabel metal2 77000 76832 77000 76832 0 net157
rlabel metal2 78176 75544 78176 75544 0 net158
rlabel metal2 73080 1134 73080 1134 0 net159
rlabel metal2 54712 74592 54712 74592 0 net16
rlabel metal2 73304 2030 73304 2030 0 net160
rlabel metal2 73528 2590 73528 2590 0 net161
rlabel metal2 30296 2030 30296 2030 0 net162
rlabel metal2 30968 2030 30968 2030 0 net163
rlabel metal2 31640 2030 31640 2030 0 net164
rlabel metal2 32312 2590 32312 2590 0 net165
rlabel metal2 32984 1246 32984 1246 0 net166
rlabel metal2 33656 2030 33656 2030 0 net167
rlabel metal2 34328 2030 34328 2030 0 net168
rlabel metal2 35000 2030 35000 2030 0 net169
rlabel metal2 51800 75992 51800 75992 0 net17
rlabel metal2 35672 2030 35672 2030 0 net170
rlabel metal2 36344 2030 36344 2030 0 net171
rlabel metal2 37016 2590 37016 2590 0 net172
rlabel metal2 37688 2030 37688 2030 0 net173
rlabel metal2 38360 2030 38360 2030 0 net174
rlabel metal2 39032 2030 39032 2030 0 net175
rlabel metal2 39704 2030 39704 2030 0 net176
rlabel metal2 40376 2030 40376 2030 0 net177
rlabel metal2 41048 2030 41048 2030 0 net178
rlabel metal2 41720 2030 41720 2030 0 net179
rlabel metal2 47320 71064 47320 71064 0 net18
rlabel metal2 42392 2030 42392 2030 0 net180
rlabel metal2 43064 2030 43064 2030 0 net181
rlabel metal2 43736 2030 43736 2030 0 net182
rlabel metal2 44408 1246 44408 1246 0 net183
rlabel metal2 45080 2030 45080 2030 0 net184
rlabel metal2 45752 1246 45752 1246 0 net185
rlabel metal2 46424 1302 46424 1302 0 net186
rlabel metal2 47096 1246 47096 1246 0 net187
rlabel metal2 47768 2030 47768 2030 0 net188
rlabel metal2 48440 1246 48440 1246 0 net189
rlabel metal2 52808 75880 52808 75880 0 net19
rlabel metal2 49112 1246 49112 1246 0 net190
rlabel metal2 49784 2030 49784 2030 0 net191
rlabel metal2 50456 1246 50456 1246 0 net192
rlabel metal2 51128 2590 51128 2590 0 net193
rlabel metal2 51800 2030 51800 2030 0 net194
rlabel metal2 52472 1246 52472 1246 0 net195
rlabel metal2 53144 2030 53144 2030 0 net196
rlabel metal2 53816 1246 53816 1246 0 net197
rlabel metal2 37128 76384 37128 76384 0 net2
rlabel metal2 62440 74928 62440 74928 0 net20
rlabel metal2 64568 74704 64568 74704 0 net21
rlabel metal2 7952 75768 7952 75768 0 net22
rlabel metal2 24808 76104 24808 76104 0 net23
rlabel metal2 26600 75040 26600 75040 0 net24
rlabel metal2 29064 75208 29064 75208 0 net25
rlabel metal2 30576 73528 30576 73528 0 net26
rlabel metal2 31528 74256 31528 74256 0 net27
rlabel metal2 32424 75432 32424 75432 0 net28
rlabel metal2 35168 75544 35168 75544 0 net29
rlabel metal2 39760 70280 39760 70280 0 net3
rlabel metal2 37128 73808 37128 73808 0 net30
rlabel metal2 12936 74088 12936 74088 0 net31
rlabel metal2 21448 73920 21448 73920 0 net32
rlabel metal2 30968 75152 30968 75152 0 net33
rlabel metal2 19880 76104 19880 76104 0 net34
rlabel metal2 20888 75880 20888 75880 0 net35
rlabel metal2 24024 75824 24024 75824 0 net36
rlabel metal2 54488 2030 54488 2030 0 net37
rlabel metal2 55160 2590 55160 2590 0 net38
rlabel metal2 55832 1246 55832 1246 0 net39
rlabel metal2 44296 70168 44296 70168 0 net4
rlabel metal2 56504 2030 56504 2030 0 net40
rlabel metal2 57176 1246 57176 1246 0 net41
rlabel metal2 57848 1302 57848 1302 0 net42
rlabel metal2 58520 2030 58520 2030 0 net43
rlabel metal2 59192 2590 59192 2590 0 net44
rlabel metal2 59864 2030 59864 2030 0 net45
rlabel metal2 60536 1246 60536 1246 0 net46
rlabel metal2 61208 1302 61208 1302 0 net47
rlabel metal2 61880 2030 61880 2030 0 net48
rlabel metal2 62552 1246 62552 1246 0 net49
rlabel metal3 44576 73528 44576 73528 0 net5
rlabel metal2 63224 2590 63224 2590 0 net50
rlabel metal2 63896 1246 63896 1246 0 net51
rlabel metal2 64568 1134 64568 1134 0 net52
rlabel metal2 65240 1134 65240 1134 0 net53
rlabel metal2 65912 1302 65912 1302 0 net54
rlabel metal2 66584 1190 66584 1190 0 net55
rlabel metal2 67256 1246 67256 1246 0 net56
rlabel metal2 67928 2030 67928 2030 0 net57
rlabel metal2 68600 1246 68600 1246 0 net58
rlabel metal2 69272 1246 69272 1246 0 net59
rlabel metal2 46760 76160 46760 76160 0 net6
rlabel metal2 69944 1302 69944 1302 0 net60
rlabel metal2 70616 2590 70616 2590 0 net61
rlabel metal2 71288 2030 71288 2030 0 net62
rlabel metal2 71960 1246 71960 1246 0 net63
rlabel metal2 72632 1246 72632 1246 0 net64
rlabel metal2 6776 2030 6776 2030 0 net65
rlabel metal2 8120 2030 8120 2030 0 net66
rlabel metal2 9016 2030 9016 2030 0 net67
rlabel metal2 9912 2030 9912 2030 0 net68
rlabel metal2 10808 2030 10808 2030 0 net69
rlabel metal2 44632 73584 44632 73584 0 net7
rlabel metal2 11704 2030 11704 2030 0 net70
rlabel metal2 12376 2030 12376 2030 0 net71
rlabel metal2 13048 2030 13048 2030 0 net72
rlabel metal2 13720 2590 13720 2590 0 net73
rlabel metal2 14392 2030 14392 2030 0 net74
rlabel metal2 15064 2030 15064 2030 0 net75
rlabel metal2 15736 2030 15736 2030 0 net76
rlabel metal2 16408 2030 16408 2030 0 net77
rlabel metal2 17080 2030 17080 2030 0 net78
rlabel metal2 17752 2590 17752 2590 0 net79
rlabel metal2 48664 72184 48664 72184 0 net8
rlabel metal2 18424 2030 18424 2030 0 net80
rlabel metal2 19096 2030 19096 2030 0 net81
rlabel metal2 19768 854 19768 854 0 net82
rlabel metal2 20440 2030 20440 2030 0 net83
rlabel metal2 21112 2030 21112 2030 0 net84
rlabel metal2 21784 2030 21784 2030 0 net85
rlabel metal2 22456 2030 22456 2030 0 net86
rlabel metal2 23128 2030 23128 2030 0 net87
rlabel metal2 23800 2030 23800 2030 0 net88
rlabel metal2 24472 2590 24472 2590 0 net89
rlabel metal2 46200 72352 46200 72352 0 net9
rlabel metal2 25144 1246 25144 1246 0 net90
rlabel metal2 25816 2030 25816 2030 0 net91
rlabel metal2 26488 2030 26488 2030 0 net92
rlabel metal2 27160 2030 27160 2030 0 net93
rlabel metal2 27832 2030 27832 2030 0 net94
rlabel metal2 28504 2030 28504 2030 0 net95
rlabel metal2 29176 2590 29176 2590 0 net96
rlabel metal2 29848 2030 29848 2030 0 net97
rlabel metal3 3416 76664 3416 76664 0 net98
rlabel metal2 4984 77938 4984 77938 0 net99
<< properties >>
string FIXED_BBOX 0 0 80000 80000
<< end >>
