magic
tech gf180mcuC
magscale 1 10
timestamp 1670287983
<< metal1 >>
rect 33842 77198 33854 77250
rect 33906 77247 33918 77250
rect 34738 77247 34750 77250
rect 33906 77201 34750 77247
rect 33906 77198 33918 77201
rect 34738 77198 34750 77201
rect 34802 77198 34814 77250
rect 42578 77086 42590 77138
rect 42642 77135 42654 77138
rect 44370 77135 44382 77138
rect 42642 77089 44382 77135
rect 42642 77086 42654 77089
rect 44370 77086 44382 77089
rect 44434 77135 44446 77138
rect 44818 77135 44830 77138
rect 44434 77089 44830 77135
rect 44434 77086 44446 77089
rect 44818 77086 44830 77089
rect 44882 77086 44894 77138
rect 40562 76974 40574 77026
rect 40626 77023 40638 77026
rect 41794 77023 41806 77026
rect 40626 76977 41806 77023
rect 40626 76974 40638 76977
rect 41794 76974 41806 76977
rect 41858 77023 41870 77026
rect 42690 77023 42702 77026
rect 41858 76977 42702 77023
rect 41858 76974 41870 76977
rect 42690 76974 42702 76977
rect 42754 76974 42766 77026
rect 46610 76974 46622 77026
rect 46674 77023 46686 77026
rect 46834 77023 46846 77026
rect 46674 76977 46846 77023
rect 46674 76974 46686 76977
rect 46834 76974 46846 76977
rect 46898 77023 46910 77026
rect 48850 77023 48862 77026
rect 46898 76977 48862 77023
rect 46898 76974 46910 76977
rect 48850 76974 48862 76977
rect 48914 76974 48926 77026
rect 60722 76974 60734 77026
rect 60786 77023 60798 77026
rect 61954 77023 61966 77026
rect 60786 76977 61966 77023
rect 60786 76974 60798 76977
rect 61954 76974 61966 76977
rect 62018 76974 62030 77026
rect 1344 76858 78624 76892
rect 1344 76806 19838 76858
rect 19890 76806 19942 76858
rect 19994 76806 20046 76858
rect 20098 76806 50558 76858
rect 50610 76806 50662 76858
rect 50714 76806 50766 76858
rect 50818 76806 78624 76858
rect 1344 76772 78624 76806
rect 5854 76690 5906 76702
rect 5854 76626 5906 76638
rect 6526 76690 6578 76702
rect 6526 76626 6578 76638
rect 7198 76690 7250 76702
rect 7198 76626 7250 76638
rect 7870 76690 7922 76702
rect 7870 76626 7922 76638
rect 9214 76690 9266 76702
rect 9214 76626 9266 76638
rect 9886 76690 9938 76702
rect 9886 76626 9938 76638
rect 11230 76690 11282 76702
rect 11230 76626 11282 76638
rect 40910 76690 40962 76702
rect 40910 76626 40962 76638
rect 43822 76690 43874 76702
rect 43822 76626 43874 76638
rect 60510 76690 60562 76702
rect 60510 76626 60562 76638
rect 61966 76690 62018 76702
rect 61966 76626 62018 76638
rect 69358 76690 69410 76702
rect 69358 76626 69410 76638
rect 69918 76690 69970 76702
rect 69918 76626 69970 76638
rect 70478 76690 70530 76702
rect 70478 76626 70530 76638
rect 70926 76690 70978 76702
rect 70926 76626 70978 76638
rect 44606 76578 44658 76590
rect 1922 76526 1934 76578
rect 1986 76526 1998 76578
rect 3938 76526 3950 76578
rect 4002 76526 4014 76578
rect 12002 76526 12014 76578
rect 12066 76526 12078 76578
rect 14018 76526 14030 76578
rect 14082 76526 14094 76578
rect 16034 76526 16046 76578
rect 16098 76526 16110 76578
rect 18050 76526 18062 76578
rect 18114 76526 18126 76578
rect 19842 76526 19854 76578
rect 19906 76526 19918 76578
rect 22082 76526 22094 76578
rect 22146 76526 22158 76578
rect 24098 76526 24110 76578
rect 24162 76526 24174 76578
rect 26114 76526 26126 76578
rect 26178 76526 26190 76578
rect 37874 76526 37886 76578
rect 37938 76526 37950 76578
rect 39106 76526 39118 76578
rect 39170 76526 39182 76578
rect 42690 76526 42702 76578
rect 42754 76526 42766 76578
rect 44606 76514 44658 76526
rect 45502 76578 45554 76590
rect 45502 76514 45554 76526
rect 45838 76578 45890 76590
rect 49870 76578 49922 76590
rect 58942 76578 58994 76590
rect 48850 76526 48862 76578
rect 48914 76526 48926 76578
rect 52882 76526 52894 76578
rect 52946 76526 52958 76578
rect 53890 76526 53902 76578
rect 53954 76526 53966 76578
rect 55010 76526 55022 76578
rect 55074 76526 55086 76578
rect 57922 76526 57934 76578
rect 57986 76526 57998 76578
rect 45838 76514 45890 76526
rect 49870 76514 49922 76526
rect 58942 76514 58994 76526
rect 59838 76578 59890 76590
rect 61618 76526 61630 76578
rect 61682 76526 61694 76578
rect 64978 76526 64990 76578
rect 65042 76526 65054 76578
rect 68002 76526 68014 76578
rect 68066 76526 68078 76578
rect 69010 76526 69022 76578
rect 69074 76526 69086 76578
rect 73042 76526 73054 76578
rect 73106 76526 73118 76578
rect 77634 76526 77646 76578
rect 77698 76526 77710 76578
rect 59838 76514 59890 76526
rect 54238 76466 54290 76478
rect 62414 76466 62466 76478
rect 5058 76414 5070 76466
rect 5122 76414 5134 76466
rect 13122 76414 13134 76466
rect 13186 76414 13198 76466
rect 15138 76414 15150 76466
rect 15202 76414 15214 76466
rect 16930 76414 16942 76466
rect 16994 76414 17006 76466
rect 19170 76414 19182 76466
rect 19234 76414 19246 76466
rect 20962 76414 20974 76466
rect 21026 76414 21038 76466
rect 23202 76414 23214 76466
rect 23266 76414 23278 76466
rect 24994 76414 25006 76466
rect 25058 76414 25070 76466
rect 27234 76414 27246 76466
rect 27298 76414 27310 76466
rect 28242 76414 28254 76466
rect 28306 76414 28318 76466
rect 30034 76414 30046 76466
rect 30098 76414 30110 76466
rect 32162 76414 32174 76466
rect 32226 76414 32238 76466
rect 34066 76414 34078 76466
rect 34130 76414 34142 76466
rect 36082 76414 36094 76466
rect 36146 76414 36158 76466
rect 38098 76414 38110 76466
rect 38162 76414 38174 76466
rect 44818 76414 44830 76466
rect 44882 76414 44894 76466
rect 50082 76414 50094 76466
rect 50146 76414 50158 76466
rect 50306 76414 50318 76466
rect 50370 76414 50382 76466
rect 59154 76414 59166 76466
rect 59218 76414 59230 76466
rect 54238 76402 54290 76414
rect 62414 76402 62466 76414
rect 46398 76354 46450 76366
rect 3266 76302 3278 76354
rect 3330 76302 3342 76354
rect 28802 76302 28814 76354
rect 28866 76302 28878 76354
rect 30706 76302 30718 76354
rect 30770 76302 30782 76354
rect 32722 76302 32734 76354
rect 32786 76302 32798 76354
rect 34738 76302 34750 76354
rect 34802 76302 34814 76354
rect 36754 76302 36766 76354
rect 36818 76302 36830 76354
rect 40002 76302 40014 76354
rect 40066 76302 40078 76354
rect 41682 76302 41694 76354
rect 41746 76302 41758 76354
rect 46398 76290 46450 76302
rect 51102 76354 51154 76366
rect 56130 76302 56142 76354
rect 56194 76302 56206 76354
rect 56914 76302 56926 76354
rect 56978 76302 56990 76354
rect 51102 76290 51154 76302
rect 43710 76242 43762 76254
rect 43710 76178 43762 76190
rect 44046 76242 44098 76254
rect 44046 76178 44098 76190
rect 46734 76242 46786 76254
rect 46734 76178 46786 76190
rect 49758 76242 49810 76254
rect 49758 76178 49810 76190
rect 62862 76242 62914 76254
rect 62862 76178 62914 76190
rect 65886 76242 65938 76254
rect 65886 76178 65938 76190
rect 74510 76242 74562 76254
rect 74510 76178 74562 76190
rect 1344 76074 78624 76108
rect 1344 76022 4478 76074
rect 4530 76022 4582 76074
rect 4634 76022 4686 76074
rect 4738 76022 35198 76074
rect 35250 76022 35302 76074
rect 35354 76022 35406 76074
rect 35458 76022 65918 76074
rect 65970 76022 66022 76074
rect 66074 76022 66126 76074
rect 66178 76022 78624 76074
rect 1344 75988 78624 76022
rect 29486 75906 29538 75918
rect 29486 75842 29538 75854
rect 44718 75906 44770 75918
rect 44718 75842 44770 75854
rect 53118 75906 53170 75918
rect 53118 75842 53170 75854
rect 1822 75794 1874 75806
rect 1822 75730 1874 75742
rect 19854 75794 19906 75806
rect 19854 75730 19906 75742
rect 20974 75794 21026 75806
rect 20974 75730 21026 75742
rect 23998 75794 24050 75806
rect 23998 75730 24050 75742
rect 26798 75794 26850 75806
rect 26798 75730 26850 75742
rect 29374 75794 29426 75806
rect 29374 75730 29426 75742
rect 35086 75794 35138 75806
rect 40462 75794 40514 75806
rect 36306 75742 36318 75794
rect 36370 75742 36382 75794
rect 38770 75742 38782 75794
rect 38834 75742 38846 75794
rect 35086 75730 35138 75742
rect 40462 75730 40514 75742
rect 44830 75794 44882 75806
rect 44830 75730 44882 75742
rect 48414 75794 48466 75806
rect 65214 75794 65266 75806
rect 48962 75742 48974 75794
rect 49026 75742 49038 75794
rect 75058 75742 75070 75794
rect 75122 75742 75134 75794
rect 48414 75730 48466 75742
rect 65214 75730 65266 75742
rect 13806 75682 13858 75694
rect 13806 75618 13858 75630
rect 15822 75682 15874 75694
rect 15822 75618 15874 75630
rect 17838 75682 17890 75694
rect 30382 75682 30434 75694
rect 30034 75630 30046 75682
rect 30098 75630 30110 75682
rect 17838 75618 17890 75630
rect 30382 75618 30434 75630
rect 30606 75682 30658 75694
rect 30606 75618 30658 75630
rect 31166 75682 31218 75694
rect 31166 75618 31218 75630
rect 31390 75682 31442 75694
rect 40686 75682 40738 75694
rect 31714 75630 31726 75682
rect 31778 75630 31790 75682
rect 38098 75630 38110 75682
rect 38162 75630 38174 75682
rect 31390 75618 31442 75630
rect 40686 75618 40738 75630
rect 41134 75682 41186 75694
rect 50430 75682 50482 75694
rect 46722 75630 46734 75682
rect 46786 75630 46798 75682
rect 49074 75630 49086 75682
rect 49138 75630 49150 75682
rect 41134 75618 41186 75630
rect 50430 75618 50482 75630
rect 52334 75682 52386 75694
rect 52334 75618 52386 75630
rect 53006 75682 53058 75694
rect 54462 75682 54514 75694
rect 54114 75630 54126 75682
rect 54178 75630 54190 75682
rect 53006 75618 53058 75630
rect 54462 75618 54514 75630
rect 55134 75682 55186 75694
rect 59614 75682 59666 75694
rect 55570 75630 55582 75682
rect 55634 75630 55646 75682
rect 55134 75618 55186 75630
rect 59614 75618 59666 75630
rect 3166 75570 3218 75582
rect 3166 75506 3218 75518
rect 5182 75570 5234 75582
rect 5182 75506 5234 75518
rect 13246 75570 13298 75582
rect 13246 75506 13298 75518
rect 15262 75570 15314 75582
rect 15262 75506 15314 75518
rect 17278 75570 17330 75582
rect 17278 75506 17330 75518
rect 19294 75570 19346 75582
rect 19294 75506 19346 75518
rect 21758 75570 21810 75582
rect 21758 75506 21810 75518
rect 23326 75570 23378 75582
rect 23326 75506 23378 75518
rect 25342 75570 25394 75582
rect 25342 75506 25394 75518
rect 27358 75570 27410 75582
rect 27358 75506 27410 75518
rect 28254 75570 28306 75582
rect 28254 75506 28306 75518
rect 28590 75570 28642 75582
rect 28590 75506 28642 75518
rect 29262 75570 29314 75582
rect 29262 75506 29314 75518
rect 32286 75570 32338 75582
rect 32286 75506 32338 75518
rect 32622 75570 32674 75582
rect 32622 75506 32674 75518
rect 33182 75570 33234 75582
rect 33182 75506 33234 75518
rect 33518 75570 33570 75582
rect 33518 75506 33570 75518
rect 33742 75570 33794 75582
rect 33742 75506 33794 75518
rect 34414 75570 34466 75582
rect 34414 75506 34466 75518
rect 34974 75570 35026 75582
rect 34974 75506 35026 75518
rect 35310 75570 35362 75582
rect 35310 75506 35362 75518
rect 35534 75570 35586 75582
rect 35534 75506 35586 75518
rect 36654 75570 36706 75582
rect 36654 75506 36706 75518
rect 36878 75570 36930 75582
rect 36878 75506 36930 75518
rect 40014 75570 40066 75582
rect 40014 75506 40066 75518
rect 41694 75570 41746 75582
rect 41694 75506 41746 75518
rect 42254 75570 42306 75582
rect 42254 75506 42306 75518
rect 42926 75570 42978 75582
rect 42926 75506 42978 75518
rect 43038 75570 43090 75582
rect 43038 75506 43090 75518
rect 43486 75570 43538 75582
rect 43486 75506 43538 75518
rect 43822 75570 43874 75582
rect 43822 75506 43874 75518
rect 45950 75570 46002 75582
rect 45950 75506 46002 75518
rect 47406 75570 47458 75582
rect 47406 75506 47458 75518
rect 49422 75570 49474 75582
rect 49422 75506 49474 75518
rect 53790 75570 53842 75582
rect 53790 75506 53842 75518
rect 56478 75570 56530 75582
rect 56478 75506 56530 75518
rect 57374 75570 57426 75582
rect 57374 75506 57426 75518
rect 59166 75570 59218 75582
rect 59166 75506 59218 75518
rect 59950 75570 60002 75582
rect 59950 75506 60002 75518
rect 60510 75570 60562 75582
rect 60510 75506 60562 75518
rect 63086 75570 63138 75582
rect 63086 75506 63138 75518
rect 63758 75570 63810 75582
rect 63758 75506 63810 75518
rect 64430 75570 64482 75582
rect 64430 75506 64482 75518
rect 65662 75570 65714 75582
rect 65662 75506 65714 75518
rect 66334 75570 66386 75582
rect 70702 75570 70754 75582
rect 69010 75518 69022 75570
rect 69074 75518 69086 75570
rect 66334 75506 66386 75518
rect 70702 75506 70754 75518
rect 71710 75570 71762 75582
rect 71710 75506 71762 75518
rect 72382 75570 72434 75582
rect 72382 75506 72434 75518
rect 73390 75570 73442 75582
rect 73390 75506 73442 75518
rect 73950 75570 74002 75582
rect 77982 75570 78034 75582
rect 76962 75518 76974 75570
rect 77026 75518 77038 75570
rect 73950 75506 74002 75518
rect 77982 75506 78034 75518
rect 33294 75458 33346 75470
rect 33294 75394 33346 75406
rect 36318 75458 36370 75470
rect 36318 75394 36370 75406
rect 36430 75458 36482 75470
rect 36430 75394 36482 75406
rect 37550 75458 37602 75470
rect 37550 75394 37602 75406
rect 40126 75458 40178 75470
rect 40126 75394 40178 75406
rect 40238 75458 40290 75470
rect 40238 75394 40290 75406
rect 41246 75458 41298 75470
rect 41246 75394 41298 75406
rect 41470 75458 41522 75470
rect 41470 75394 41522 75406
rect 42478 75458 42530 75470
rect 42478 75394 42530 75406
rect 42702 75458 42754 75470
rect 42702 75394 42754 75406
rect 43710 75458 43762 75470
rect 43710 75394 43762 75406
rect 43934 75458 43986 75470
rect 43934 75394 43986 75406
rect 44046 75458 44098 75470
rect 44046 75394 44098 75406
rect 44942 75458 44994 75470
rect 44942 75394 44994 75406
rect 45614 75458 45666 75470
rect 45614 75394 45666 75406
rect 46510 75458 46562 75470
rect 48302 75458 48354 75470
rect 47730 75406 47742 75458
rect 47794 75406 47806 75458
rect 46510 75394 46562 75406
rect 48302 75394 48354 75406
rect 49534 75458 49586 75470
rect 49534 75394 49586 75406
rect 49758 75458 49810 75470
rect 49758 75394 49810 75406
rect 50878 75458 50930 75470
rect 50878 75394 50930 75406
rect 50990 75458 51042 75470
rect 50990 75394 51042 75406
rect 51102 75458 51154 75470
rect 51102 75394 51154 75406
rect 51662 75458 51714 75470
rect 51662 75394 51714 75406
rect 51774 75458 51826 75470
rect 51774 75394 51826 75406
rect 51886 75458 51938 75470
rect 51886 75394 51938 75406
rect 52894 75458 52946 75470
rect 52894 75394 52946 75406
rect 53902 75458 53954 75470
rect 53902 75394 53954 75406
rect 54014 75458 54066 75470
rect 54014 75394 54066 75406
rect 55022 75458 55074 75470
rect 55022 75394 55074 75406
rect 55246 75458 55298 75470
rect 55246 75394 55298 75406
rect 56142 75458 56194 75470
rect 56142 75394 56194 75406
rect 57038 75458 57090 75470
rect 58270 75458 58322 75470
rect 57922 75406 57934 75458
rect 57986 75406 57998 75458
rect 57038 75394 57090 75406
rect 58270 75394 58322 75406
rect 58830 75458 58882 75470
rect 58830 75394 58882 75406
rect 59838 75458 59890 75470
rect 59838 75394 59890 75406
rect 61742 75458 61794 75470
rect 61742 75394 61794 75406
rect 62414 75458 62466 75470
rect 62414 75394 62466 75406
rect 66894 75458 66946 75470
rect 66894 75394 66946 75406
rect 70030 75458 70082 75470
rect 70030 75394 70082 75406
rect 73054 75458 73106 75470
rect 73054 75394 73106 75406
rect 1344 75290 78624 75324
rect 1344 75238 19838 75290
rect 19890 75238 19942 75290
rect 19994 75238 20046 75290
rect 20098 75238 50558 75290
rect 50610 75238 50662 75290
rect 50714 75238 50766 75290
rect 50818 75238 78624 75290
rect 1344 75204 78624 75238
rect 28702 75122 28754 75134
rect 28702 75058 28754 75070
rect 29374 75122 29426 75134
rect 29374 75058 29426 75070
rect 30270 75122 30322 75134
rect 30270 75058 30322 75070
rect 31278 75122 31330 75134
rect 34638 75122 34690 75134
rect 33170 75070 33182 75122
rect 33234 75070 33246 75122
rect 31278 75058 31330 75070
rect 34638 75058 34690 75070
rect 35646 75122 35698 75134
rect 35646 75058 35698 75070
rect 35758 75122 35810 75134
rect 35758 75058 35810 75070
rect 36430 75122 36482 75134
rect 36430 75058 36482 75070
rect 38782 75122 38834 75134
rect 38782 75058 38834 75070
rect 40014 75122 40066 75134
rect 40014 75058 40066 75070
rect 40126 75122 40178 75134
rect 40126 75058 40178 75070
rect 41022 75122 41074 75134
rect 44942 75122 44994 75134
rect 43138 75070 43150 75122
rect 43202 75070 43214 75122
rect 41022 75058 41074 75070
rect 44942 75058 44994 75070
rect 45950 75122 46002 75134
rect 45950 75058 46002 75070
rect 47070 75122 47122 75134
rect 47070 75058 47122 75070
rect 54350 75122 54402 75134
rect 54350 75058 54402 75070
rect 54798 75122 54850 75134
rect 54798 75058 54850 75070
rect 56590 75122 56642 75134
rect 56590 75058 56642 75070
rect 59278 75122 59330 75134
rect 59278 75058 59330 75070
rect 62190 75122 62242 75134
rect 62190 75058 62242 75070
rect 62862 75122 62914 75134
rect 62862 75058 62914 75070
rect 63870 75122 63922 75134
rect 63870 75058 63922 75070
rect 66782 75122 66834 75134
rect 66782 75058 66834 75070
rect 67678 75122 67730 75134
rect 67678 75058 67730 75070
rect 70814 75122 70866 75134
rect 70814 75058 70866 75070
rect 72830 75122 72882 75134
rect 72830 75058 72882 75070
rect 74398 75122 74450 75134
rect 74398 75058 74450 75070
rect 75742 75122 75794 75134
rect 75742 75058 75794 75070
rect 76414 75122 76466 75134
rect 76414 75058 76466 75070
rect 77422 75122 77474 75134
rect 77422 75058 77474 75070
rect 78094 75122 78146 75134
rect 78094 75058 78146 75070
rect 29934 75010 29986 75022
rect 29934 74946 29986 74958
rect 30830 75010 30882 75022
rect 38670 75010 38722 75022
rect 37314 74958 37326 75010
rect 37378 74958 37390 75010
rect 30830 74946 30882 74958
rect 38670 74946 38722 74958
rect 39006 75010 39058 75022
rect 39006 74946 39058 74958
rect 43710 75010 43762 75022
rect 43710 74946 43762 74958
rect 47182 75010 47234 75022
rect 49982 75010 50034 75022
rect 48850 74958 48862 75010
rect 48914 74958 48926 75010
rect 49074 74958 49086 75010
rect 49138 74958 49150 75010
rect 47182 74946 47234 74958
rect 49982 74946 50034 74958
rect 52670 75010 52722 75022
rect 52670 74946 52722 74958
rect 53006 75010 53058 75022
rect 53006 74946 53058 74958
rect 53566 75010 53618 75022
rect 60174 75010 60226 75022
rect 57474 74958 57486 75010
rect 57538 74958 57550 75010
rect 53566 74946 53618 74958
rect 60174 74946 60226 74958
rect 61630 75010 61682 75022
rect 61630 74946 61682 74958
rect 31054 74898 31106 74910
rect 31054 74834 31106 74846
rect 31390 74898 31442 74910
rect 31390 74834 31442 74846
rect 32062 74898 32114 74910
rect 32062 74834 32114 74846
rect 33742 74898 33794 74910
rect 35534 74898 35586 74910
rect 39454 74898 39506 74910
rect 34402 74846 34414 74898
rect 34466 74846 34478 74898
rect 35186 74846 35198 74898
rect 35250 74846 35262 74898
rect 37538 74846 37550 74898
rect 37602 74846 37614 74898
rect 38210 74846 38222 74898
rect 38274 74846 38286 74898
rect 33742 74834 33794 74846
rect 35534 74834 35586 74846
rect 39454 74834 39506 74846
rect 39902 74898 39954 74910
rect 42478 74898 42530 74910
rect 40786 74846 40798 74898
rect 40850 74846 40862 74898
rect 39902 74834 39954 74846
rect 42478 74834 42530 74846
rect 42590 74898 42642 74910
rect 42590 74834 42642 74846
rect 42702 74898 42754 74910
rect 44158 74898 44210 74910
rect 45726 74898 45778 74910
rect 43922 74846 43934 74898
rect 43986 74846 43998 74898
rect 44482 74846 44494 74898
rect 44546 74846 44558 74898
rect 42702 74834 42754 74846
rect 44158 74834 44210 74846
rect 45726 74834 45778 74846
rect 46846 74898 46898 74910
rect 46846 74834 46898 74846
rect 50318 74898 50370 74910
rect 54014 74898 54066 74910
rect 58830 74898 58882 74910
rect 59502 74898 59554 74910
rect 51426 74846 51438 74898
rect 51490 74846 51502 74898
rect 53778 74846 53790 74898
rect 53842 74846 53854 74898
rect 54338 74846 54350 74898
rect 54402 74846 54414 74898
rect 57698 74846 57710 74898
rect 57762 74846 57774 74898
rect 59154 74846 59166 74898
rect 59218 74846 59230 74898
rect 50318 74834 50370 74846
rect 54014 74834 54066 74846
rect 58830 74834 58882 74846
rect 59502 74834 59554 74846
rect 61518 74898 61570 74910
rect 61518 74834 61570 74846
rect 29262 74786 29314 74798
rect 29262 74722 29314 74734
rect 32286 74786 32338 74798
rect 41694 74786 41746 74798
rect 38658 74734 38670 74786
rect 38722 74734 38734 74786
rect 32286 74722 32338 74734
rect 41694 74722 41746 74734
rect 43822 74786 43874 74798
rect 43822 74722 43874 74734
rect 45838 74786 45890 74798
rect 45838 74722 45890 74734
rect 46174 74786 46226 74798
rect 46174 74722 46226 74734
rect 50990 74786 51042 74798
rect 55694 74786 55746 74798
rect 51874 74734 51886 74786
rect 51938 74734 51950 74786
rect 50990 74722 51042 74734
rect 55694 74722 55746 74734
rect 58270 74786 58322 74798
rect 58270 74722 58322 74734
rect 59390 74786 59442 74798
rect 59390 74722 59442 74734
rect 60286 74786 60338 74798
rect 60286 74722 60338 74734
rect 60958 74786 61010 74798
rect 60958 74722 61010 74734
rect 63422 74786 63474 74798
rect 63422 74722 63474 74734
rect 33518 74674 33570 74686
rect 32610 74622 32622 74674
rect 32674 74622 32686 74674
rect 33518 74610 33570 74622
rect 36766 74674 36818 74686
rect 46398 74674 46450 74686
rect 44594 74622 44606 74674
rect 44658 74671 44670 74674
rect 44930 74671 44942 74674
rect 44658 74625 44942 74671
rect 44658 74622 44670 74625
rect 44930 74622 44942 74625
rect 44994 74622 45006 74674
rect 36766 74610 36818 74622
rect 46398 74610 46450 74622
rect 48190 74674 48242 74686
rect 48190 74610 48242 74622
rect 48526 74674 48578 74686
rect 48526 74610 48578 74622
rect 55246 74674 55298 74686
rect 55246 74610 55298 74622
rect 55470 74674 55522 74686
rect 55470 74610 55522 74622
rect 56926 74674 56978 74686
rect 56926 74610 56978 74622
rect 60846 74674 60898 74686
rect 60846 74610 60898 74622
rect 1344 74506 78624 74540
rect 1344 74454 4478 74506
rect 4530 74454 4582 74506
rect 4634 74454 4686 74506
rect 4738 74454 35198 74506
rect 35250 74454 35302 74506
rect 35354 74454 35406 74506
rect 35458 74454 65918 74506
rect 65970 74454 66022 74506
rect 66074 74454 66126 74506
rect 66178 74454 78624 74506
rect 1344 74420 78624 74454
rect 34302 74338 34354 74350
rect 35422 74338 35474 74350
rect 33954 74286 33966 74338
rect 34018 74286 34030 74338
rect 35074 74286 35086 74338
rect 35138 74286 35150 74338
rect 34302 74274 34354 74286
rect 35422 74274 35474 74286
rect 36318 74338 36370 74350
rect 36318 74274 36370 74286
rect 38222 74338 38274 74350
rect 38222 74274 38274 74286
rect 44270 74338 44322 74350
rect 44270 74274 44322 74286
rect 48638 74338 48690 74350
rect 50766 74338 50818 74350
rect 49298 74286 49310 74338
rect 49362 74286 49374 74338
rect 48638 74274 48690 74286
rect 50766 74274 50818 74286
rect 28926 74226 28978 74238
rect 28926 74162 28978 74174
rect 29262 74226 29314 74238
rect 29262 74162 29314 74174
rect 29822 74226 29874 74238
rect 29822 74162 29874 74174
rect 34526 74226 34578 74238
rect 34526 74162 34578 74174
rect 35646 74226 35698 74238
rect 35646 74162 35698 74174
rect 40462 74226 40514 74238
rect 43934 74226 43986 74238
rect 42018 74174 42030 74226
rect 42082 74174 42094 74226
rect 40462 74162 40514 74174
rect 43934 74162 43986 74174
rect 44830 74226 44882 74238
rect 44830 74162 44882 74174
rect 47854 74226 47906 74238
rect 61630 74226 61682 74238
rect 53218 74174 53230 74226
rect 53282 74174 53294 74226
rect 47854 74162 47906 74174
rect 61630 74162 61682 74174
rect 62526 74226 62578 74238
rect 62526 74162 62578 74174
rect 62974 74226 63026 74238
rect 62974 74162 63026 74174
rect 63534 74226 63586 74238
rect 63534 74162 63586 74174
rect 78094 74226 78146 74238
rect 78094 74162 78146 74174
rect 31166 74114 31218 74126
rect 30482 74062 30494 74114
rect 30546 74062 30558 74114
rect 31166 74050 31218 74062
rect 32062 74114 32114 74126
rect 32062 74050 32114 74062
rect 33070 74114 33122 74126
rect 33070 74050 33122 74062
rect 36654 74114 36706 74126
rect 38110 74114 38162 74126
rect 37426 74062 37438 74114
rect 37490 74062 37502 74114
rect 36654 74050 36706 74062
rect 38110 74050 38162 74062
rect 38782 74114 38834 74126
rect 40350 74114 40402 74126
rect 44158 74114 44210 74126
rect 39330 74062 39342 74114
rect 39394 74062 39406 74114
rect 41682 74062 41694 74114
rect 41746 74062 41758 74114
rect 42914 74062 42926 74114
rect 42978 74062 42990 74114
rect 43138 74062 43150 74114
rect 43202 74062 43214 74114
rect 38782 74050 38834 74062
rect 40350 74050 40402 74062
rect 44158 74050 44210 74062
rect 45502 74114 45554 74126
rect 48750 74114 48802 74126
rect 50654 74114 50706 74126
rect 46050 74062 46062 74114
rect 46114 74062 46126 74114
rect 50082 74062 50094 74114
rect 50146 74062 50158 74114
rect 45502 74050 45554 74062
rect 48750 74050 48802 74062
rect 50654 74050 50706 74062
rect 51326 74114 51378 74126
rect 51326 74050 51378 74062
rect 52110 74114 52162 74126
rect 54686 74114 54738 74126
rect 52882 74062 52894 74114
rect 52946 74062 52958 74114
rect 53890 74062 53902 74114
rect 53954 74062 53966 74114
rect 54226 74062 54238 74114
rect 54290 74062 54302 74114
rect 52110 74050 52162 74062
rect 54686 74050 54738 74062
rect 55022 74114 55074 74126
rect 55022 74050 55074 74062
rect 55694 74114 55746 74126
rect 55694 74050 55746 74062
rect 57598 74114 57650 74126
rect 57598 74050 57650 74062
rect 58718 74114 58770 74126
rect 58718 74050 58770 74062
rect 58942 74114 58994 74126
rect 62078 74114 62130 74126
rect 59266 74062 59278 74114
rect 59330 74062 59342 74114
rect 58942 74050 58994 74062
rect 62078 74050 62130 74062
rect 32398 74002 32450 74014
rect 39902 74002 39954 74014
rect 37202 73950 37214 74002
rect 37266 73950 37278 74002
rect 32398 73938 32450 73950
rect 39902 73938 39954 73950
rect 40574 74002 40626 74014
rect 40574 73938 40626 73950
rect 40798 74002 40850 74014
rect 45614 74002 45666 74014
rect 42130 73950 42142 74002
rect 42194 73950 42206 74002
rect 40798 73938 40850 73950
rect 45614 73938 45666 73950
rect 45726 74002 45778 74014
rect 45726 73938 45778 73950
rect 49758 74002 49810 74014
rect 49758 73938 49810 73950
rect 49870 74002 49922 74014
rect 49870 73938 49922 73950
rect 50878 74002 50930 74014
rect 50878 73938 50930 73950
rect 51102 74002 51154 74014
rect 51102 73938 51154 73950
rect 51998 74002 52050 74014
rect 56030 74002 56082 74014
rect 52770 73950 52782 74002
rect 52834 73950 52846 74002
rect 51998 73938 52050 73950
rect 56030 73938 56082 73950
rect 56814 74002 56866 74014
rect 56814 73938 56866 73950
rect 57038 74002 57090 74014
rect 57038 73938 57090 73950
rect 57934 74002 57986 74014
rect 57934 73938 57986 73950
rect 30270 73890 30322 73902
rect 30270 73826 30322 73838
rect 31502 73890 31554 73902
rect 31502 73826 31554 73838
rect 33406 73890 33458 73902
rect 33406 73826 33458 73838
rect 38894 73890 38946 73902
rect 38894 73826 38946 73838
rect 39006 73890 39058 73902
rect 39006 73826 39058 73838
rect 44270 73890 44322 73902
rect 44270 73826 44322 73838
rect 46622 73890 46674 73902
rect 46622 73826 46674 73838
rect 47294 73890 47346 73902
rect 47294 73826 47346 73838
rect 48638 73890 48690 73902
rect 48638 73826 48690 73838
rect 51774 73890 51826 73902
rect 51774 73826 51826 73838
rect 54910 73890 54962 73902
rect 54910 73826 54962 73838
rect 55806 73890 55858 73902
rect 55806 73826 55858 73838
rect 56926 73890 56978 73902
rect 56926 73826 56978 73838
rect 57822 73890 57874 73902
rect 57822 73826 57874 73838
rect 58830 73890 58882 73902
rect 58830 73826 58882 73838
rect 59838 73890 59890 73902
rect 59838 73826 59890 73838
rect 60510 73890 60562 73902
rect 60510 73826 60562 73838
rect 1344 73722 78624 73756
rect 1344 73670 19838 73722
rect 19890 73670 19942 73722
rect 19994 73670 20046 73722
rect 20098 73670 50558 73722
rect 50610 73670 50662 73722
rect 50714 73670 50766 73722
rect 50818 73670 78624 73722
rect 1344 73636 78624 73670
rect 30942 73554 30994 73566
rect 30942 73490 30994 73502
rect 31390 73554 31442 73566
rect 31390 73490 31442 73502
rect 32174 73554 32226 73566
rect 32174 73490 32226 73502
rect 32734 73554 32786 73566
rect 32734 73490 32786 73502
rect 33406 73554 33458 73566
rect 33406 73490 33458 73502
rect 33518 73554 33570 73566
rect 33518 73490 33570 73502
rect 34526 73554 34578 73566
rect 34526 73490 34578 73502
rect 35422 73554 35474 73566
rect 35422 73490 35474 73502
rect 36318 73554 36370 73566
rect 36318 73490 36370 73502
rect 36654 73554 36706 73566
rect 36654 73490 36706 73502
rect 36878 73554 36930 73566
rect 36878 73490 36930 73502
rect 39678 73554 39730 73566
rect 39678 73490 39730 73502
rect 40910 73554 40962 73566
rect 40910 73490 40962 73502
rect 42254 73554 42306 73566
rect 42254 73490 42306 73502
rect 47854 73554 47906 73566
rect 47854 73490 47906 73502
rect 48526 73554 48578 73566
rect 48526 73490 48578 73502
rect 50318 73554 50370 73566
rect 50318 73490 50370 73502
rect 54574 73554 54626 73566
rect 54574 73490 54626 73502
rect 55358 73554 55410 73566
rect 55358 73490 55410 73502
rect 55918 73554 55970 73566
rect 55918 73490 55970 73502
rect 56030 73554 56082 73566
rect 56030 73490 56082 73502
rect 60398 73554 60450 73566
rect 60398 73490 60450 73502
rect 60958 73554 61010 73566
rect 60958 73490 61010 73502
rect 61406 73554 61458 73566
rect 61406 73490 61458 73502
rect 61854 73554 61906 73566
rect 61854 73490 61906 73502
rect 33630 73442 33682 73454
rect 33630 73378 33682 73390
rect 34190 73442 34242 73454
rect 34190 73378 34242 73390
rect 35310 73442 35362 73454
rect 35310 73378 35362 73390
rect 35982 73442 36034 73454
rect 35982 73378 36034 73390
rect 36094 73442 36146 73454
rect 36094 73378 36146 73390
rect 37550 73442 37602 73454
rect 37550 73378 37602 73390
rect 37886 73442 37938 73454
rect 37886 73378 37938 73390
rect 40574 73442 40626 73454
rect 40574 73378 40626 73390
rect 44606 73442 44658 73454
rect 44606 73378 44658 73390
rect 44718 73442 44770 73454
rect 44718 73378 44770 73390
rect 47182 73442 47234 73454
rect 47182 73378 47234 73390
rect 50878 73442 50930 73454
rect 50878 73378 50930 73390
rect 51102 73442 51154 73454
rect 51102 73378 51154 73390
rect 52894 73442 52946 73454
rect 52894 73378 52946 73390
rect 54014 73442 54066 73454
rect 54014 73378 54066 73390
rect 54910 73442 54962 73454
rect 54910 73378 54962 73390
rect 57262 73442 57314 73454
rect 57262 73378 57314 73390
rect 36990 73330 37042 73342
rect 36990 73266 37042 73278
rect 38446 73330 38498 73342
rect 38446 73266 38498 73278
rect 40798 73330 40850 73342
rect 40798 73266 40850 73278
rect 41022 73330 41074 73342
rect 41022 73266 41074 73278
rect 43150 73330 43202 73342
rect 43150 73266 43202 73278
rect 44158 73330 44210 73342
rect 44158 73266 44210 73278
rect 44382 73330 44434 73342
rect 47294 73330 47346 73342
rect 53566 73330 53618 73342
rect 45938 73278 45950 73330
rect 46002 73278 46014 73330
rect 51202 73278 51214 73330
rect 51266 73327 51278 73330
rect 51538 73327 51550 73330
rect 51266 73281 51550 73327
rect 51266 73278 51278 73281
rect 51538 73278 51550 73281
rect 51602 73278 51614 73330
rect 52434 73278 52446 73330
rect 52498 73278 52510 73330
rect 44382 73266 44434 73278
rect 47294 73266 47346 73278
rect 53566 73266 53618 73278
rect 53678 73330 53730 73342
rect 53678 73266 53730 73278
rect 53902 73330 53954 73342
rect 53902 73266 53954 73278
rect 56142 73330 56194 73342
rect 56142 73266 56194 73278
rect 56590 73330 56642 73342
rect 57698 73278 57710 73330
rect 57762 73278 57774 73330
rect 59266 73278 59278 73330
rect 59330 73278 59342 73330
rect 56590 73266 56642 73278
rect 30382 73218 30434 73230
rect 30382 73154 30434 73166
rect 39790 73218 39842 73230
rect 39790 73154 39842 73166
rect 41694 73218 41746 73230
rect 41694 73154 41746 73166
rect 42702 73218 42754 73230
rect 42702 73154 42754 73166
rect 45502 73218 45554 73230
rect 47966 73218 48018 73230
rect 45826 73166 45838 73218
rect 45890 73166 45902 73218
rect 45502 73154 45554 73166
rect 47966 73154 48018 73166
rect 49422 73218 49474 73230
rect 58830 73218 58882 73230
rect 50754 73166 50766 73218
rect 50818 73166 50830 73218
rect 52098 73166 52110 73218
rect 52162 73166 52174 73218
rect 58034 73166 58046 73218
rect 58098 73166 58110 73218
rect 59602 73166 59614 73218
rect 59666 73166 59678 73218
rect 49422 73154 49474 73166
rect 58830 73154 58882 73166
rect 38670 73106 38722 73118
rect 39902 73106 39954 73118
rect 38994 73054 39006 73106
rect 39058 73054 39070 73106
rect 38670 73042 38722 73054
rect 39902 73042 39954 73054
rect 42926 73106 42978 73118
rect 42926 73042 42978 73054
rect 44942 73106 44994 73118
rect 44942 73042 44994 73054
rect 47182 73106 47234 73118
rect 47182 73042 47234 73054
rect 49646 73106 49698 73118
rect 49646 73042 49698 73054
rect 49870 73106 49922 73118
rect 49870 73042 49922 73054
rect 1344 72938 78624 72972
rect 1344 72886 4478 72938
rect 4530 72886 4582 72938
rect 4634 72886 4686 72938
rect 4738 72886 35198 72938
rect 35250 72886 35302 72938
rect 35354 72886 35406 72938
rect 35458 72886 65918 72938
rect 65970 72886 66022 72938
rect 66074 72886 66126 72938
rect 66178 72886 78624 72938
rect 1344 72852 78624 72886
rect 55582 72770 55634 72782
rect 33730 72718 33742 72770
rect 33794 72767 33806 72770
rect 34290 72767 34302 72770
rect 33794 72721 34302 72767
rect 33794 72718 33806 72721
rect 34290 72718 34302 72721
rect 34354 72718 34366 72770
rect 57138 72718 57150 72770
rect 57202 72718 57214 72770
rect 55582 72706 55634 72718
rect 31950 72658 32002 72670
rect 31950 72594 32002 72606
rect 32398 72658 32450 72670
rect 32398 72594 32450 72606
rect 32846 72658 32898 72670
rect 32846 72594 32898 72606
rect 33294 72658 33346 72670
rect 33294 72594 33346 72606
rect 33742 72658 33794 72670
rect 33742 72594 33794 72606
rect 34190 72658 34242 72670
rect 34190 72594 34242 72606
rect 35422 72658 35474 72670
rect 35422 72594 35474 72606
rect 36990 72658 37042 72670
rect 49758 72658 49810 72670
rect 43138 72606 43150 72658
rect 43202 72606 43214 72658
rect 43922 72606 43934 72658
rect 43986 72606 43998 72658
rect 45602 72606 45614 72658
rect 45666 72606 45678 72658
rect 36990 72594 37042 72606
rect 49758 72594 49810 72606
rect 50878 72658 50930 72670
rect 54910 72658 54962 72670
rect 59278 72658 59330 72670
rect 51538 72606 51550 72658
rect 51602 72606 51614 72658
rect 56466 72606 56478 72658
rect 56530 72606 56542 72658
rect 58034 72606 58046 72658
rect 58098 72606 58110 72658
rect 50878 72594 50930 72606
rect 54910 72594 54962 72606
rect 59278 72594 59330 72606
rect 59726 72658 59778 72670
rect 59726 72594 59778 72606
rect 60174 72658 60226 72670
rect 60174 72594 60226 72606
rect 60622 72658 60674 72670
rect 60622 72594 60674 72606
rect 37886 72546 37938 72558
rect 37426 72494 37438 72546
rect 37490 72494 37502 72546
rect 37886 72482 37938 72494
rect 39006 72546 39058 72558
rect 40350 72546 40402 72558
rect 46286 72546 46338 72558
rect 39666 72494 39678 72546
rect 39730 72494 39742 72546
rect 39890 72494 39902 72546
rect 39954 72494 39966 72546
rect 40562 72494 40574 72546
rect 40626 72494 40638 72546
rect 42802 72494 42814 72546
rect 42866 72494 42878 72546
rect 45154 72494 45166 72546
rect 45218 72494 45230 72546
rect 39006 72482 39058 72494
rect 40350 72482 40402 72494
rect 46286 72482 46338 72494
rect 46622 72546 46674 72558
rect 46622 72482 46674 72494
rect 49646 72546 49698 72558
rect 49646 72482 49698 72494
rect 49870 72546 49922 72558
rect 49870 72482 49922 72494
rect 50766 72546 50818 72558
rect 54686 72546 54738 72558
rect 51874 72494 51886 72546
rect 51938 72494 51950 72546
rect 52434 72494 52446 72546
rect 52498 72494 52510 72546
rect 53330 72494 53342 72546
rect 53394 72494 53406 72546
rect 50766 72482 50818 72494
rect 54686 72482 54738 72494
rect 55694 72546 55746 72558
rect 57026 72494 57038 72546
rect 57090 72494 57102 72546
rect 57250 72494 57262 72546
rect 57314 72494 57326 72546
rect 57922 72494 57934 72546
rect 57986 72494 57998 72546
rect 55694 72482 55746 72494
rect 34750 72434 34802 72446
rect 34750 72370 34802 72382
rect 36430 72434 36482 72446
rect 36430 72370 36482 72382
rect 40238 72434 40290 72446
rect 40238 72370 40290 72382
rect 42254 72434 42306 72446
rect 42254 72370 42306 72382
rect 43934 72434 43986 72446
rect 43934 72370 43986 72382
rect 44158 72434 44210 72446
rect 44158 72370 44210 72382
rect 44718 72434 44770 72446
rect 44718 72370 44770 72382
rect 46398 72434 46450 72446
rect 46398 72370 46450 72382
rect 47070 72434 47122 72446
rect 47070 72370 47122 72382
rect 48190 72434 48242 72446
rect 48190 72370 48242 72382
rect 49086 72434 49138 72446
rect 49086 72370 49138 72382
rect 50094 72434 50146 72446
rect 55582 72434 55634 72446
rect 51650 72382 51662 72434
rect 51714 72382 51726 72434
rect 52658 72382 52670 72434
rect 52722 72382 52734 72434
rect 54338 72382 54350 72434
rect 54402 72382 54414 72434
rect 50094 72370 50146 72382
rect 55582 72370 55634 72382
rect 59166 72434 59218 72446
rect 59166 72370 59218 72382
rect 35310 72322 35362 72334
rect 35310 72258 35362 72270
rect 38558 72322 38610 72334
rect 38558 72258 38610 72270
rect 41694 72322 41746 72334
rect 41694 72258 41746 72270
rect 47630 72322 47682 72334
rect 47630 72258 47682 72270
rect 1344 72154 78624 72188
rect 1344 72102 19838 72154
rect 19890 72102 19942 72154
rect 19994 72102 20046 72154
rect 20098 72102 50558 72154
rect 50610 72102 50662 72154
rect 50714 72102 50766 72154
rect 50818 72102 78624 72154
rect 1344 72068 78624 72102
rect 33854 71986 33906 71998
rect 33854 71922 33906 71934
rect 35982 71986 36034 71998
rect 35982 71922 36034 71934
rect 36430 71986 36482 71998
rect 36430 71922 36482 71934
rect 36990 71986 37042 71998
rect 36990 71922 37042 71934
rect 37438 71986 37490 71998
rect 37438 71922 37490 71934
rect 37662 71986 37714 71998
rect 41022 71986 41074 71998
rect 45726 71986 45778 71998
rect 38434 71934 38446 71986
rect 38498 71934 38510 71986
rect 43026 71934 43038 71986
rect 43090 71934 43102 71986
rect 37662 71922 37714 71934
rect 41022 71922 41074 71934
rect 45726 71922 45778 71934
rect 47182 71986 47234 71998
rect 47182 71922 47234 71934
rect 47630 71986 47682 71998
rect 47630 71922 47682 71934
rect 48078 71986 48130 71998
rect 48078 71922 48130 71934
rect 52334 71986 52386 71998
rect 52334 71922 52386 71934
rect 54462 71986 54514 71998
rect 58718 71986 58770 71998
rect 58034 71934 58046 71986
rect 58098 71934 58110 71986
rect 54462 71922 54514 71934
rect 58718 71922 58770 71934
rect 59278 71986 59330 71998
rect 59278 71922 59330 71934
rect 59614 71986 59666 71998
rect 59614 71922 59666 71934
rect 37774 71874 37826 71886
rect 45166 71874 45218 71886
rect 40114 71822 40126 71874
rect 40178 71822 40190 71874
rect 43250 71822 43262 71874
rect 43314 71822 43326 71874
rect 43922 71822 43934 71874
rect 43986 71822 43998 71874
rect 37774 71810 37826 71822
rect 45166 71810 45218 71822
rect 49422 71874 49474 71886
rect 49422 71810 49474 71822
rect 53006 71874 53058 71886
rect 53006 71810 53058 71822
rect 55470 71874 55522 71886
rect 56690 71822 56702 71874
rect 56754 71822 56766 71874
rect 57922 71822 57934 71874
rect 57986 71822 57998 71874
rect 55470 71810 55522 71822
rect 44494 71762 44546 71774
rect 38994 71710 39006 71762
rect 39058 71710 39070 71762
rect 39778 71710 39790 71762
rect 39842 71710 39854 71762
rect 41794 71710 41806 71762
rect 41858 71710 41870 71762
rect 42802 71710 42814 71762
rect 42866 71710 42878 71762
rect 43586 71710 43598 71762
rect 43650 71710 43662 71762
rect 44494 71698 44546 71710
rect 44942 71762 44994 71774
rect 45938 71710 45950 71762
rect 46002 71759 46014 71762
rect 46162 71759 46174 71762
rect 46002 71713 46174 71759
rect 46002 71710 46014 71713
rect 46162 71710 46174 71713
rect 46226 71710 46238 71762
rect 50194 71710 50206 71762
rect 50258 71710 50270 71762
rect 51538 71710 51550 71762
rect 51602 71710 51614 71762
rect 53218 71710 53230 71762
rect 53282 71710 53294 71762
rect 53554 71710 53566 71762
rect 53618 71710 53630 71762
rect 55234 71710 55246 71762
rect 55298 71710 55310 71762
rect 56914 71710 56926 71762
rect 56978 71710 56990 71762
rect 44942 71698 44994 71710
rect 34974 71650 35026 71662
rect 34974 71586 35026 71598
rect 35422 71650 35474 71662
rect 35422 71586 35474 71598
rect 44718 71650 44770 71662
rect 44718 71586 44770 71598
rect 46286 71650 46338 71662
rect 46286 71586 46338 71598
rect 46734 71650 46786 71662
rect 46734 71586 46786 71598
rect 48526 71650 48578 71662
rect 51650 71598 51662 71650
rect 51714 71598 51726 71650
rect 48526 71586 48578 71598
rect 34862 71538 34914 71550
rect 46050 71486 46062 71538
rect 46114 71535 46126 71538
rect 46722 71535 46734 71538
rect 46114 71489 46734 71535
rect 46114 71486 46126 71489
rect 46722 71486 46734 71489
rect 46786 71486 46798 71538
rect 47954 71486 47966 71538
rect 48018 71535 48030 71538
rect 48514 71535 48526 71538
rect 48018 71489 48526 71535
rect 48018 71486 48030 71489
rect 48514 71486 48526 71489
rect 48578 71486 48590 71538
rect 34862 71474 34914 71486
rect 1344 71370 78624 71404
rect 1344 71318 4478 71370
rect 4530 71318 4582 71370
rect 4634 71318 4686 71370
rect 4738 71318 35198 71370
rect 35250 71318 35302 71370
rect 35354 71318 35406 71370
rect 35458 71318 65918 71370
rect 65970 71318 66022 71370
rect 66074 71318 66126 71370
rect 66178 71318 78624 71370
rect 1344 71284 78624 71318
rect 39902 71202 39954 71214
rect 56142 71202 56194 71214
rect 57374 71202 57426 71214
rect 41570 71150 41582 71202
rect 41634 71150 41646 71202
rect 45602 71150 45614 71202
rect 45666 71199 45678 71202
rect 46274 71199 46286 71202
rect 45666 71153 46286 71199
rect 45666 71150 45678 71153
rect 46274 71150 46286 71153
rect 46338 71150 46350 71202
rect 46498 71150 46510 71202
rect 46562 71199 46574 71202
rect 46946 71199 46958 71202
rect 46562 71153 46958 71199
rect 46562 71150 46574 71153
rect 46946 71150 46958 71153
rect 47010 71150 47022 71202
rect 54450 71150 54462 71202
rect 54514 71199 54526 71202
rect 54674 71199 54686 71202
rect 54514 71153 54686 71199
rect 54514 71150 54526 71153
rect 54674 71150 54686 71153
rect 54738 71199 54750 71202
rect 54898 71199 54910 71202
rect 54738 71153 54910 71199
rect 54738 71150 54750 71153
rect 54898 71150 54910 71153
rect 54962 71150 54974 71202
rect 56466 71150 56478 71202
rect 56530 71150 56542 71202
rect 39902 71138 39954 71150
rect 56142 71138 56194 71150
rect 57374 71138 57426 71150
rect 35198 71090 35250 71102
rect 35198 71026 35250 71038
rect 35646 71090 35698 71102
rect 35646 71026 35698 71038
rect 37326 71090 37378 71102
rect 37326 71026 37378 71038
rect 37662 71090 37714 71102
rect 37662 71026 37714 71038
rect 38222 71090 38274 71102
rect 42142 71090 42194 71102
rect 40898 71038 40910 71090
rect 40962 71038 40974 71090
rect 38222 71026 38274 71038
rect 42142 71026 42194 71038
rect 45614 71090 45666 71102
rect 45614 71026 45666 71038
rect 46062 71090 46114 71102
rect 46062 71026 46114 71038
rect 46958 71090 47010 71102
rect 46958 71026 47010 71038
rect 47406 71090 47458 71102
rect 47406 71026 47458 71038
rect 47854 71090 47906 71102
rect 47854 71026 47906 71038
rect 48750 71090 48802 71102
rect 48750 71026 48802 71038
rect 49310 71090 49362 71102
rect 49310 71026 49362 71038
rect 50878 71090 50930 71102
rect 50878 71026 50930 71038
rect 51326 71090 51378 71102
rect 51326 71026 51378 71038
rect 51886 71090 51938 71102
rect 51886 71026 51938 71038
rect 52894 71090 52946 71102
rect 52894 71026 52946 71038
rect 53230 71090 53282 71102
rect 53230 71026 53282 71038
rect 54126 71090 54178 71102
rect 54126 71026 54178 71038
rect 54462 71090 54514 71102
rect 54462 71026 54514 71038
rect 54910 71090 54962 71102
rect 54910 71026 54962 71038
rect 57262 71090 57314 71102
rect 57262 71026 57314 71038
rect 57934 71090 57986 71102
rect 57934 71026 57986 71038
rect 36430 70978 36482 70990
rect 36430 70914 36482 70926
rect 39006 70978 39058 70990
rect 42814 70978 42866 70990
rect 44270 70978 44322 70990
rect 46510 70978 46562 70990
rect 41122 70926 41134 70978
rect 41186 70926 41198 70978
rect 43586 70926 43598 70978
rect 43650 70926 43662 70978
rect 44930 70926 44942 70978
rect 44994 70926 45006 70978
rect 39006 70914 39058 70926
rect 42814 70914 42866 70926
rect 44270 70914 44322 70926
rect 46510 70914 46562 70926
rect 51774 70978 51826 70990
rect 51774 70914 51826 70926
rect 52110 70978 52162 70990
rect 52110 70914 52162 70926
rect 52334 70978 52386 70990
rect 52334 70914 52386 70926
rect 55918 70978 55970 70990
rect 57026 70926 57038 70978
rect 57090 70926 57102 70978
rect 55918 70914 55970 70926
rect 38670 70866 38722 70878
rect 38670 70802 38722 70814
rect 39790 70866 39842 70878
rect 39790 70802 39842 70814
rect 50206 70866 50258 70878
rect 50206 70802 50258 70814
rect 36094 70754 36146 70766
rect 36094 70690 36146 70702
rect 39902 70754 39954 70766
rect 39902 70690 39954 70702
rect 48302 70754 48354 70766
rect 48302 70690 48354 70702
rect 49646 70754 49698 70766
rect 49646 70690 49698 70702
rect 55470 70754 55522 70766
rect 55470 70690 55522 70702
rect 1344 70586 78624 70620
rect 1344 70534 19838 70586
rect 19890 70534 19942 70586
rect 19994 70534 20046 70586
rect 20098 70534 50558 70586
rect 50610 70534 50662 70586
rect 50714 70534 50766 70586
rect 50818 70534 78624 70586
rect 1344 70500 78624 70534
rect 38110 70418 38162 70430
rect 38110 70354 38162 70366
rect 38558 70418 38610 70430
rect 38558 70354 38610 70366
rect 39006 70418 39058 70430
rect 39006 70354 39058 70366
rect 39454 70418 39506 70430
rect 39454 70354 39506 70366
rect 40126 70418 40178 70430
rect 40126 70354 40178 70366
rect 40350 70418 40402 70430
rect 40350 70354 40402 70366
rect 41022 70418 41074 70430
rect 43934 70418 43986 70430
rect 42802 70366 42814 70418
rect 42866 70366 42878 70418
rect 41022 70354 41074 70366
rect 43934 70354 43986 70366
rect 44270 70418 44322 70430
rect 44270 70354 44322 70366
rect 44830 70418 44882 70430
rect 44830 70354 44882 70366
rect 45278 70418 45330 70430
rect 45278 70354 45330 70366
rect 45726 70418 45778 70430
rect 45726 70354 45778 70366
rect 46174 70418 46226 70430
rect 46174 70354 46226 70366
rect 46622 70418 46674 70430
rect 46622 70354 46674 70366
rect 47182 70418 47234 70430
rect 47182 70354 47234 70366
rect 49758 70418 49810 70430
rect 49758 70354 49810 70366
rect 50206 70418 50258 70430
rect 50206 70354 50258 70366
rect 50654 70418 50706 70430
rect 50654 70354 50706 70366
rect 51102 70418 51154 70430
rect 51102 70354 51154 70366
rect 51662 70418 51714 70430
rect 51662 70354 51714 70366
rect 52558 70418 52610 70430
rect 52558 70354 52610 70366
rect 53006 70418 53058 70430
rect 53006 70354 53058 70366
rect 54238 70418 54290 70430
rect 54238 70354 54290 70366
rect 54686 70418 54738 70430
rect 54686 70354 54738 70366
rect 55358 70418 55410 70430
rect 55358 70354 55410 70366
rect 56030 70418 56082 70430
rect 56030 70354 56082 70366
rect 56478 70418 56530 70430
rect 56478 70354 56530 70366
rect 40462 70306 40514 70318
rect 40462 70242 40514 70254
rect 56926 70306 56978 70318
rect 56926 70242 56978 70254
rect 37214 70194 37266 70206
rect 37214 70130 37266 70142
rect 37550 70194 37602 70206
rect 37550 70130 37602 70142
rect 43150 70194 43202 70206
rect 43150 70130 43202 70142
rect 43374 70194 43426 70206
rect 43374 70130 43426 70142
rect 39566 70082 39618 70094
rect 39566 70018 39618 70030
rect 53454 70082 53506 70094
rect 53454 70018 53506 70030
rect 37986 69918 37998 69970
rect 38050 69967 38062 69970
rect 38546 69967 38558 69970
rect 38050 69921 38558 69967
rect 38050 69918 38062 69921
rect 38546 69918 38558 69921
rect 38610 69918 38622 69970
rect 43698 69918 43710 69970
rect 43762 69967 43774 69970
rect 44706 69967 44718 69970
rect 43762 69921 44718 69967
rect 43762 69918 43774 69921
rect 44706 69918 44718 69921
rect 44770 69918 44782 69970
rect 1344 69802 78624 69836
rect 1344 69750 4478 69802
rect 4530 69750 4582 69802
rect 4634 69750 4686 69802
rect 4738 69750 35198 69802
rect 35250 69750 35302 69802
rect 35354 69750 35406 69802
rect 35458 69750 65918 69802
rect 65970 69750 66022 69802
rect 66074 69750 66126 69802
rect 66178 69750 78624 69802
rect 1344 69716 78624 69750
rect 38558 69522 38610 69534
rect 38558 69458 38610 69470
rect 39006 69522 39058 69534
rect 39006 69458 39058 69470
rect 39678 69522 39730 69534
rect 39678 69458 39730 69470
rect 40126 69522 40178 69534
rect 40126 69458 40178 69470
rect 43262 69522 43314 69534
rect 43262 69458 43314 69470
rect 44494 69522 44546 69534
rect 44494 69458 44546 69470
rect 44830 69522 44882 69534
rect 44830 69458 44882 69470
rect 54686 69522 54738 69534
rect 54686 69458 54738 69470
rect 1344 69018 78624 69052
rect 1344 68966 19838 69018
rect 19890 68966 19942 69018
rect 19994 68966 20046 69018
rect 20098 68966 50558 69018
rect 50610 68966 50662 69018
rect 50714 68966 50766 69018
rect 50818 68966 78624 69018
rect 1344 68932 78624 68966
rect 1344 68234 78624 68268
rect 1344 68182 4478 68234
rect 4530 68182 4582 68234
rect 4634 68182 4686 68234
rect 4738 68182 35198 68234
rect 35250 68182 35302 68234
rect 35354 68182 35406 68234
rect 35458 68182 65918 68234
rect 65970 68182 66022 68234
rect 66074 68182 66126 68234
rect 66178 68182 78624 68234
rect 1344 68148 78624 68182
rect 1344 67450 78624 67484
rect 1344 67398 19838 67450
rect 19890 67398 19942 67450
rect 19994 67398 20046 67450
rect 20098 67398 50558 67450
rect 50610 67398 50662 67450
rect 50714 67398 50766 67450
rect 50818 67398 78624 67450
rect 1344 67364 78624 67398
rect 1344 66666 78624 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 35198 66666
rect 35250 66614 35302 66666
rect 35354 66614 35406 66666
rect 35458 66614 65918 66666
rect 65970 66614 66022 66666
rect 66074 66614 66126 66666
rect 66178 66614 78624 66666
rect 1344 66580 78624 66614
rect 1344 65882 78624 65916
rect 1344 65830 19838 65882
rect 19890 65830 19942 65882
rect 19994 65830 20046 65882
rect 20098 65830 50558 65882
rect 50610 65830 50662 65882
rect 50714 65830 50766 65882
rect 50818 65830 78624 65882
rect 1344 65796 78624 65830
rect 1344 65098 78624 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 35198 65098
rect 35250 65046 35302 65098
rect 35354 65046 35406 65098
rect 35458 65046 65918 65098
rect 65970 65046 66022 65098
rect 66074 65046 66126 65098
rect 66178 65046 78624 65098
rect 1344 65012 78624 65046
rect 1344 64314 78624 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 50558 64314
rect 50610 64262 50662 64314
rect 50714 64262 50766 64314
rect 50818 64262 78624 64314
rect 1344 64228 78624 64262
rect 1344 63530 78624 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 65918 63530
rect 65970 63478 66022 63530
rect 66074 63478 66126 63530
rect 66178 63478 78624 63530
rect 1344 63444 78624 63478
rect 1344 62746 78624 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 50558 62746
rect 50610 62694 50662 62746
rect 50714 62694 50766 62746
rect 50818 62694 78624 62746
rect 1344 62660 78624 62694
rect 1344 61962 78624 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 65918 61962
rect 65970 61910 66022 61962
rect 66074 61910 66126 61962
rect 66178 61910 78624 61962
rect 1344 61876 78624 61910
rect 1344 61178 78624 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 50558 61178
rect 50610 61126 50662 61178
rect 50714 61126 50766 61178
rect 50818 61126 78624 61178
rect 1344 61092 78624 61126
rect 1344 60394 78624 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 65918 60394
rect 65970 60342 66022 60394
rect 66074 60342 66126 60394
rect 66178 60342 78624 60394
rect 1344 60308 78624 60342
rect 1344 59610 78624 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 50558 59610
rect 50610 59558 50662 59610
rect 50714 59558 50766 59610
rect 50818 59558 78624 59610
rect 1344 59524 78624 59558
rect 1344 58826 78624 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 65918 58826
rect 65970 58774 66022 58826
rect 66074 58774 66126 58826
rect 66178 58774 78624 58826
rect 1344 58740 78624 58774
rect 1344 58042 78624 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 50558 58042
rect 50610 57990 50662 58042
rect 50714 57990 50766 58042
rect 50818 57990 78624 58042
rect 1344 57956 78624 57990
rect 1344 57258 78624 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 65918 57258
rect 65970 57206 66022 57258
rect 66074 57206 66126 57258
rect 66178 57206 78624 57258
rect 1344 57172 78624 57206
rect 1344 56474 78624 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 78624 56474
rect 1344 56388 78624 56422
rect 1344 55690 78624 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 65918 55690
rect 65970 55638 66022 55690
rect 66074 55638 66126 55690
rect 66178 55638 78624 55690
rect 1344 55604 78624 55638
rect 1344 54906 78624 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 78624 54906
rect 1344 54820 78624 54854
rect 1344 54122 78624 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 65918 54122
rect 65970 54070 66022 54122
rect 66074 54070 66126 54122
rect 66178 54070 78624 54122
rect 1344 54036 78624 54070
rect 1344 53338 78624 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 78624 53338
rect 1344 53252 78624 53286
rect 1344 52554 78624 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 65918 52554
rect 65970 52502 66022 52554
rect 66074 52502 66126 52554
rect 66178 52502 78624 52554
rect 1344 52468 78624 52502
rect 1344 51770 78624 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 78624 51770
rect 1344 51684 78624 51718
rect 1344 50986 78624 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 65918 50986
rect 65970 50934 66022 50986
rect 66074 50934 66126 50986
rect 66178 50934 78624 50986
rect 1344 50900 78624 50934
rect 1344 50202 78624 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 78624 50202
rect 1344 50116 78624 50150
rect 1344 49418 78624 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 65918 49418
rect 65970 49366 66022 49418
rect 66074 49366 66126 49418
rect 66178 49366 78624 49418
rect 1344 49332 78624 49366
rect 1344 48634 78624 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 78624 48634
rect 1344 48548 78624 48582
rect 1344 47850 78624 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 65918 47850
rect 65970 47798 66022 47850
rect 66074 47798 66126 47850
rect 66178 47798 78624 47850
rect 1344 47764 78624 47798
rect 1344 47066 78624 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 78624 47066
rect 1344 46980 78624 47014
rect 1344 46282 78624 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 65918 46282
rect 65970 46230 66022 46282
rect 66074 46230 66126 46282
rect 66178 46230 78624 46282
rect 1344 46196 78624 46230
rect 1344 45498 78624 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 78624 45498
rect 1344 45412 78624 45446
rect 1344 44714 78624 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 65918 44714
rect 65970 44662 66022 44714
rect 66074 44662 66126 44714
rect 66178 44662 78624 44714
rect 1344 44628 78624 44662
rect 1344 43930 78624 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 78624 43930
rect 1344 43844 78624 43878
rect 1344 43146 78624 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 65918 43146
rect 65970 43094 66022 43146
rect 66074 43094 66126 43146
rect 66178 43094 78624 43146
rect 1344 43060 78624 43094
rect 1344 42362 78624 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 78624 42362
rect 1344 42276 78624 42310
rect 1344 41578 78624 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 65918 41578
rect 65970 41526 66022 41578
rect 66074 41526 66126 41578
rect 66178 41526 78624 41578
rect 1344 41492 78624 41526
rect 1344 40794 78624 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 78624 40794
rect 1344 40708 78624 40742
rect 1344 40010 78624 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 65918 40010
rect 65970 39958 66022 40010
rect 66074 39958 66126 40010
rect 66178 39958 78624 40010
rect 1344 39924 78624 39958
rect 1344 39226 78624 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 78624 39226
rect 1344 39140 78624 39174
rect 1344 38442 78624 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 65918 38442
rect 65970 38390 66022 38442
rect 66074 38390 66126 38442
rect 66178 38390 78624 38442
rect 1344 38356 78624 38390
rect 1344 37658 78624 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 78624 37658
rect 1344 37572 78624 37606
rect 1344 36874 78624 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 65918 36874
rect 65970 36822 66022 36874
rect 66074 36822 66126 36874
rect 66178 36822 78624 36874
rect 1344 36788 78624 36822
rect 1344 36090 78624 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 78624 36090
rect 1344 36004 78624 36038
rect 1344 35306 78624 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 65918 35306
rect 65970 35254 66022 35306
rect 66074 35254 66126 35306
rect 66178 35254 78624 35306
rect 1344 35220 78624 35254
rect 1344 34522 78624 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 78624 34522
rect 1344 34436 78624 34470
rect 1344 33738 78624 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 65918 33738
rect 65970 33686 66022 33738
rect 66074 33686 66126 33738
rect 66178 33686 78624 33738
rect 1344 33652 78624 33686
rect 1344 32954 78624 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 78624 32954
rect 1344 32868 78624 32902
rect 1344 32170 78624 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 65918 32170
rect 65970 32118 66022 32170
rect 66074 32118 66126 32170
rect 66178 32118 78624 32170
rect 1344 32084 78624 32118
rect 1344 31386 78624 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 78624 31386
rect 1344 31300 78624 31334
rect 1344 30602 78624 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 65918 30602
rect 65970 30550 66022 30602
rect 66074 30550 66126 30602
rect 66178 30550 78624 30602
rect 1344 30516 78624 30550
rect 1344 29818 78624 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 78624 29818
rect 1344 29732 78624 29766
rect 1344 29034 78624 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 65918 29034
rect 65970 28982 66022 29034
rect 66074 28982 66126 29034
rect 66178 28982 78624 29034
rect 1344 28948 78624 28982
rect 1344 28250 78624 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 78624 28250
rect 1344 28164 78624 28198
rect 1344 27466 78624 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 65918 27466
rect 65970 27414 66022 27466
rect 66074 27414 66126 27466
rect 66178 27414 78624 27466
rect 1344 27380 78624 27414
rect 1344 26682 78624 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 78624 26682
rect 1344 26596 78624 26630
rect 1344 25898 78624 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 65918 25898
rect 65970 25846 66022 25898
rect 66074 25846 66126 25898
rect 66178 25846 78624 25898
rect 1344 25812 78624 25846
rect 1344 25114 78624 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 78624 25114
rect 1344 25028 78624 25062
rect 1344 24330 78624 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 65918 24330
rect 65970 24278 66022 24330
rect 66074 24278 66126 24330
rect 66178 24278 78624 24330
rect 1344 24244 78624 24278
rect 1344 23546 78624 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 78624 23546
rect 1344 23460 78624 23494
rect 1344 22762 78624 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 65918 22762
rect 65970 22710 66022 22762
rect 66074 22710 66126 22762
rect 66178 22710 78624 22762
rect 1344 22676 78624 22710
rect 1344 21978 78624 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 78624 21978
rect 1344 21892 78624 21926
rect 1344 21194 78624 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 65918 21194
rect 65970 21142 66022 21194
rect 66074 21142 66126 21194
rect 66178 21142 78624 21194
rect 1344 21108 78624 21142
rect 1344 20410 78624 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 78624 20410
rect 1344 20324 78624 20358
rect 1344 19626 78624 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 65918 19626
rect 65970 19574 66022 19626
rect 66074 19574 66126 19626
rect 66178 19574 78624 19626
rect 1344 19540 78624 19574
rect 1344 18842 78624 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 78624 18842
rect 1344 18756 78624 18790
rect 1344 18058 78624 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 65918 18058
rect 65970 18006 66022 18058
rect 66074 18006 66126 18058
rect 66178 18006 78624 18058
rect 1344 17972 78624 18006
rect 1344 17274 78624 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 78624 17274
rect 1344 17188 78624 17222
rect 1344 16490 78624 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 65918 16490
rect 65970 16438 66022 16490
rect 66074 16438 66126 16490
rect 66178 16438 78624 16490
rect 1344 16404 78624 16438
rect 1344 15706 78624 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 78624 15706
rect 1344 15620 78624 15654
rect 1344 14922 78624 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 65918 14922
rect 65970 14870 66022 14922
rect 66074 14870 66126 14922
rect 66178 14870 78624 14922
rect 1344 14836 78624 14870
rect 1344 14138 78624 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 78624 14138
rect 1344 14052 78624 14086
rect 1344 13354 78624 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 65918 13354
rect 65970 13302 66022 13354
rect 66074 13302 66126 13354
rect 66178 13302 78624 13354
rect 1344 13268 78624 13302
rect 1344 12570 78624 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 78624 12570
rect 1344 12484 78624 12518
rect 1344 11786 78624 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 65918 11786
rect 65970 11734 66022 11786
rect 66074 11734 66126 11786
rect 66178 11734 78624 11786
rect 1344 11700 78624 11734
rect 1344 11002 78624 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 78624 11002
rect 1344 10916 78624 10950
rect 1344 10218 78624 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 65918 10218
rect 65970 10166 66022 10218
rect 66074 10166 66126 10218
rect 66178 10166 78624 10218
rect 1344 10132 78624 10166
rect 1344 9434 78624 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 78624 9434
rect 1344 9348 78624 9382
rect 1344 8650 78624 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 65918 8650
rect 65970 8598 66022 8650
rect 66074 8598 66126 8650
rect 66178 8598 78624 8650
rect 1344 8564 78624 8598
rect 1344 7866 78624 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 78624 7866
rect 1344 7780 78624 7814
rect 1344 7082 78624 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 65918 7082
rect 65970 7030 66022 7082
rect 66074 7030 66126 7082
rect 66178 7030 78624 7082
rect 1344 6996 78624 7030
rect 1344 6298 78624 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 78624 6298
rect 1344 6212 78624 6246
rect 1344 5514 78624 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 65918 5514
rect 65970 5462 66022 5514
rect 66074 5462 66126 5514
rect 66178 5462 78624 5514
rect 1344 5428 78624 5462
rect 1344 4730 78624 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 78624 4730
rect 1344 4644 78624 4678
rect 73278 4450 73330 4462
rect 73278 4386 73330 4398
rect 73950 4450 74002 4462
rect 73950 4386 74002 4398
rect 1344 3946 78624 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 65918 3946
rect 65970 3894 66022 3946
rect 66074 3894 66126 3946
rect 66178 3894 78624 3946
rect 1344 3860 78624 3894
rect 6974 3330 7026 3342
rect 6974 3266 7026 3278
rect 8318 3330 8370 3342
rect 8318 3266 8370 3278
rect 9214 3330 9266 3342
rect 9214 3266 9266 3278
rect 10110 3330 10162 3342
rect 10110 3266 10162 3278
rect 10782 3330 10834 3342
rect 10782 3266 10834 3278
rect 11566 3330 11618 3342
rect 11566 3266 11618 3278
rect 12238 3330 12290 3342
rect 12238 3266 12290 3278
rect 12910 3330 12962 3342
rect 12910 3266 12962 3278
rect 13582 3330 13634 3342
rect 13582 3266 13634 3278
rect 14254 3330 14306 3342
rect 14254 3266 14306 3278
rect 14926 3330 14978 3342
rect 14926 3266 14978 3278
rect 15598 3330 15650 3342
rect 15598 3266 15650 3278
rect 16270 3330 16322 3342
rect 16270 3266 16322 3278
rect 16942 3330 16994 3342
rect 16942 3266 16994 3278
rect 17614 3330 17666 3342
rect 17614 3266 17666 3278
rect 18286 3330 18338 3342
rect 18286 3266 18338 3278
rect 18958 3330 19010 3342
rect 18958 3266 19010 3278
rect 19630 3330 19682 3342
rect 19630 3266 19682 3278
rect 20302 3330 20354 3342
rect 20302 3266 20354 3278
rect 20974 3330 21026 3342
rect 20974 3266 21026 3278
rect 21758 3330 21810 3342
rect 21758 3266 21810 3278
rect 22430 3330 22482 3342
rect 22430 3266 22482 3278
rect 23102 3330 23154 3342
rect 23102 3266 23154 3278
rect 23774 3330 23826 3342
rect 23774 3266 23826 3278
rect 24446 3330 24498 3342
rect 24446 3266 24498 3278
rect 25118 3330 25170 3342
rect 25118 3266 25170 3278
rect 25790 3330 25842 3342
rect 25790 3266 25842 3278
rect 26462 3330 26514 3342
rect 26462 3266 26514 3278
rect 27134 3330 27186 3342
rect 27134 3266 27186 3278
rect 27806 3330 27858 3342
rect 27806 3266 27858 3278
rect 28478 3330 28530 3342
rect 28478 3266 28530 3278
rect 29150 3330 29202 3342
rect 29150 3266 29202 3278
rect 29822 3330 29874 3342
rect 29822 3266 29874 3278
rect 30494 3330 30546 3342
rect 30494 3266 30546 3278
rect 31166 3330 31218 3342
rect 31166 3266 31218 3278
rect 31838 3330 31890 3342
rect 31838 3266 31890 3278
rect 32510 3330 32562 3342
rect 32510 3266 32562 3278
rect 33182 3330 33234 3342
rect 33182 3266 33234 3278
rect 33854 3330 33906 3342
rect 33854 3266 33906 3278
rect 34526 3330 34578 3342
rect 34526 3266 34578 3278
rect 35198 3330 35250 3342
rect 35198 3266 35250 3278
rect 35870 3330 35922 3342
rect 35870 3266 35922 3278
rect 36542 3330 36594 3342
rect 36542 3266 36594 3278
rect 37214 3330 37266 3342
rect 37214 3266 37266 3278
rect 37886 3330 37938 3342
rect 37886 3266 37938 3278
rect 38558 3330 38610 3342
rect 38558 3266 38610 3278
rect 39230 3330 39282 3342
rect 39230 3266 39282 3278
rect 39902 3330 39954 3342
rect 39902 3266 39954 3278
rect 40574 3330 40626 3342
rect 40574 3266 40626 3278
rect 41694 3330 41746 3342
rect 41694 3266 41746 3278
rect 42366 3330 42418 3342
rect 42366 3266 42418 3278
rect 43038 3330 43090 3342
rect 43038 3266 43090 3278
rect 43710 3330 43762 3342
rect 43710 3266 43762 3278
rect 44382 3330 44434 3342
rect 44382 3266 44434 3278
rect 45054 3330 45106 3342
rect 45054 3266 45106 3278
rect 45726 3330 45778 3342
rect 45726 3266 45778 3278
rect 46398 3330 46450 3342
rect 46398 3266 46450 3278
rect 47070 3330 47122 3342
rect 47070 3266 47122 3278
rect 47742 3330 47794 3342
rect 47742 3266 47794 3278
rect 48414 3330 48466 3342
rect 48414 3266 48466 3278
rect 49086 3330 49138 3342
rect 49086 3266 49138 3278
rect 49758 3330 49810 3342
rect 49758 3266 49810 3278
rect 50430 3330 50482 3342
rect 50430 3266 50482 3278
rect 51102 3330 51154 3342
rect 51102 3266 51154 3278
rect 51774 3330 51826 3342
rect 51774 3266 51826 3278
rect 52446 3330 52498 3342
rect 52446 3266 52498 3278
rect 53118 3330 53170 3342
rect 53118 3266 53170 3278
rect 53790 3330 53842 3342
rect 53790 3266 53842 3278
rect 54462 3330 54514 3342
rect 54462 3266 54514 3278
rect 55134 3330 55186 3342
rect 55134 3266 55186 3278
rect 55806 3330 55858 3342
rect 55806 3266 55858 3278
rect 56478 3330 56530 3342
rect 56478 3266 56530 3278
rect 57150 3330 57202 3342
rect 57150 3266 57202 3278
rect 57822 3330 57874 3342
rect 57822 3266 57874 3278
rect 58494 3330 58546 3342
rect 58494 3266 58546 3278
rect 59166 3330 59218 3342
rect 59166 3266 59218 3278
rect 59838 3330 59890 3342
rect 59838 3266 59890 3278
rect 60510 3330 60562 3342
rect 60510 3266 60562 3278
rect 61630 3330 61682 3342
rect 61630 3266 61682 3278
rect 62302 3330 62354 3342
rect 62302 3266 62354 3278
rect 62974 3330 63026 3342
rect 62974 3266 63026 3278
rect 63646 3330 63698 3342
rect 63646 3266 63698 3278
rect 64318 3330 64370 3342
rect 64318 3266 64370 3278
rect 64990 3330 65042 3342
rect 64990 3266 65042 3278
rect 65662 3330 65714 3342
rect 65662 3266 65714 3278
rect 66334 3330 66386 3342
rect 66334 3266 66386 3278
rect 67006 3330 67058 3342
rect 67006 3266 67058 3278
rect 67678 3330 67730 3342
rect 67678 3266 67730 3278
rect 68350 3330 68402 3342
rect 68350 3266 68402 3278
rect 69022 3330 69074 3342
rect 69022 3266 69074 3278
rect 69694 3330 69746 3342
rect 69694 3266 69746 3278
rect 70366 3330 70418 3342
rect 70366 3266 70418 3278
rect 71038 3330 71090 3342
rect 71038 3266 71090 3278
rect 71710 3330 71762 3342
rect 71710 3266 71762 3278
rect 72382 3330 72434 3342
rect 72382 3266 72434 3278
rect 73054 3330 73106 3342
rect 73054 3266 73106 3278
rect 73726 3330 73778 3342
rect 73726 3266 73778 3278
rect 74398 3330 74450 3342
rect 74398 3266 74450 3278
rect 1344 3162 78624 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 78624 3162
rect 1344 3076 78624 3110
rect 54562 1934 54574 1986
rect 54626 1983 54638 1986
rect 55122 1983 55134 1986
rect 54626 1937 55134 1983
rect 54626 1934 54638 1937
rect 55122 1934 55134 1937
rect 55186 1934 55198 1986
rect 42354 1822 42366 1874
rect 42418 1871 42430 1874
rect 43026 1871 43038 1874
rect 42418 1825 43038 1871
rect 42418 1822 42430 1825
rect 43026 1822 43038 1825
rect 43090 1822 43102 1874
rect 44482 1822 44494 1874
rect 44546 1871 44558 1874
rect 45042 1871 45054 1874
rect 44546 1825 45054 1871
rect 44546 1822 44558 1825
rect 45042 1822 45054 1825
rect 45106 1822 45118 1874
rect 47842 1822 47854 1874
rect 47906 1871 47918 1874
rect 48402 1871 48414 1874
rect 47906 1825 48414 1871
rect 47906 1822 47918 1825
rect 48402 1822 48414 1825
rect 48466 1822 48478 1874
rect 51202 1822 51214 1874
rect 51266 1871 51278 1874
rect 51762 1871 51774 1874
rect 51266 1825 51774 1871
rect 51266 1822 51278 1825
rect 51762 1822 51774 1825
rect 51826 1822 51838 1874
rect 57922 1822 57934 1874
rect 57986 1871 57998 1874
rect 58482 1871 58494 1874
rect 57986 1825 58494 1871
rect 57986 1822 57998 1825
rect 58482 1822 58494 1825
rect 58546 1822 58558 1874
rect 41010 1710 41022 1762
rect 41074 1759 41086 1762
rect 41682 1759 41694 1762
rect 41074 1713 41694 1759
rect 41074 1710 41086 1713
rect 41682 1710 41694 1713
rect 41746 1710 41758 1762
rect 43698 1710 43710 1762
rect 43762 1759 43774 1762
rect 44370 1759 44382 1762
rect 43762 1713 44382 1759
rect 43762 1710 43774 1713
rect 44370 1710 44382 1713
rect 44434 1710 44446 1762
rect 45714 1710 45726 1762
rect 45778 1759 45790 1762
rect 46386 1759 46398 1762
rect 45778 1713 46398 1759
rect 45778 1710 45790 1713
rect 46386 1710 46398 1713
rect 46450 1710 46462 1762
rect 47058 1710 47070 1762
rect 47122 1759 47134 1762
rect 47730 1759 47742 1762
rect 47122 1713 47742 1759
rect 47122 1710 47134 1713
rect 47730 1710 47742 1713
rect 47794 1710 47806 1762
rect 49074 1710 49086 1762
rect 49138 1759 49150 1762
rect 49746 1759 49758 1762
rect 49138 1713 49758 1759
rect 49138 1710 49150 1713
rect 49746 1710 49758 1713
rect 49810 1710 49822 1762
rect 50418 1710 50430 1762
rect 50482 1759 50494 1762
rect 51090 1759 51102 1762
rect 50482 1713 51102 1759
rect 50482 1710 50494 1713
rect 51090 1710 51102 1713
rect 51154 1710 51166 1762
rect 52434 1710 52446 1762
rect 52498 1759 52510 1762
rect 53106 1759 53118 1762
rect 52498 1713 53118 1759
rect 52498 1710 52510 1713
rect 53106 1710 53118 1713
rect 53170 1710 53182 1762
rect 53778 1710 53790 1762
rect 53842 1759 53854 1762
rect 54450 1759 54462 1762
rect 53842 1713 54462 1759
rect 53842 1710 53854 1713
rect 54450 1710 54462 1713
rect 54514 1710 54526 1762
rect 55906 1710 55918 1762
rect 55970 1759 55982 1762
rect 56466 1759 56478 1762
rect 55970 1713 56478 1759
rect 55970 1710 55982 1713
rect 56466 1710 56478 1713
rect 56530 1710 56542 1762
rect 57138 1710 57150 1762
rect 57202 1759 57214 1762
rect 57810 1759 57822 1762
rect 57202 1713 57822 1759
rect 57202 1710 57214 1713
rect 57810 1710 57822 1713
rect 57874 1710 57886 1762
rect 59154 1710 59166 1762
rect 59218 1759 59230 1762
rect 59826 1759 59838 1762
rect 59218 1713 59838 1759
rect 59218 1710 59230 1713
rect 59826 1710 59838 1713
rect 59890 1710 59902 1762
rect 60498 1710 60510 1762
rect 60562 1759 60574 1762
rect 61618 1759 61630 1762
rect 60562 1713 61630 1759
rect 60562 1710 60574 1713
rect 61618 1710 61630 1713
rect 61682 1710 61694 1762
rect 62514 1710 62526 1762
rect 62578 1759 62590 1762
rect 63634 1759 63646 1762
rect 62578 1713 63646 1759
rect 62578 1710 62590 1713
rect 63634 1710 63646 1713
rect 63698 1710 63710 1762
rect 63858 1710 63870 1762
rect 63922 1759 63934 1762
rect 64978 1759 64990 1762
rect 63922 1713 64990 1759
rect 63922 1710 63934 1713
rect 64978 1710 64990 1713
rect 65042 1710 65054 1762
rect 65874 1710 65886 1762
rect 65938 1759 65950 1762
rect 66994 1759 67006 1762
rect 65938 1713 67006 1759
rect 65938 1710 65950 1713
rect 66994 1710 67006 1713
rect 67058 1710 67070 1762
rect 67218 1710 67230 1762
rect 67282 1759 67294 1762
rect 68338 1759 68350 1762
rect 67282 1713 68350 1759
rect 67282 1710 67294 1713
rect 68338 1710 68350 1713
rect 68402 1710 68414 1762
rect 69234 1710 69246 1762
rect 69298 1759 69310 1762
rect 70354 1759 70366 1762
rect 69298 1713 70366 1759
rect 69298 1710 69310 1713
rect 70354 1710 70366 1713
rect 70418 1710 70430 1762
rect 70578 1710 70590 1762
rect 70642 1759 70654 1762
rect 71698 1759 71710 1762
rect 70642 1713 71710 1759
rect 70642 1710 70654 1713
rect 71698 1710 71710 1713
rect 71762 1710 71774 1762
rect 72594 1710 72606 1762
rect 72658 1759 72670 1762
rect 73714 1759 73726 1762
rect 72658 1713 73726 1759
rect 72658 1710 72670 1713
rect 73714 1710 73726 1713
rect 73778 1710 73790 1762
<< via1 >>
rect 33854 77198 33906 77250
rect 34750 77198 34802 77250
rect 42590 77086 42642 77138
rect 44382 77086 44434 77138
rect 44830 77086 44882 77138
rect 40574 76974 40626 77026
rect 41806 76974 41858 77026
rect 42702 76974 42754 77026
rect 46622 76974 46674 77026
rect 46846 76974 46898 77026
rect 48862 76974 48914 77026
rect 60734 76974 60786 77026
rect 61966 76974 62018 77026
rect 19838 76806 19890 76858
rect 19942 76806 19994 76858
rect 20046 76806 20098 76858
rect 50558 76806 50610 76858
rect 50662 76806 50714 76858
rect 50766 76806 50818 76858
rect 5854 76638 5906 76690
rect 6526 76638 6578 76690
rect 7198 76638 7250 76690
rect 7870 76638 7922 76690
rect 9214 76638 9266 76690
rect 9886 76638 9938 76690
rect 11230 76638 11282 76690
rect 40910 76638 40962 76690
rect 43822 76638 43874 76690
rect 60510 76638 60562 76690
rect 61966 76638 62018 76690
rect 69358 76638 69410 76690
rect 69918 76638 69970 76690
rect 70478 76638 70530 76690
rect 70926 76638 70978 76690
rect 1934 76526 1986 76578
rect 3950 76526 4002 76578
rect 12014 76526 12066 76578
rect 14030 76526 14082 76578
rect 16046 76526 16098 76578
rect 18062 76526 18114 76578
rect 19854 76526 19906 76578
rect 22094 76526 22146 76578
rect 24110 76526 24162 76578
rect 26126 76526 26178 76578
rect 37886 76526 37938 76578
rect 39118 76526 39170 76578
rect 42702 76526 42754 76578
rect 44606 76526 44658 76578
rect 45502 76526 45554 76578
rect 45838 76526 45890 76578
rect 48862 76526 48914 76578
rect 49870 76526 49922 76578
rect 52894 76526 52946 76578
rect 53902 76526 53954 76578
rect 55022 76526 55074 76578
rect 57934 76526 57986 76578
rect 58942 76526 58994 76578
rect 59838 76526 59890 76578
rect 61630 76526 61682 76578
rect 64990 76526 65042 76578
rect 68014 76526 68066 76578
rect 69022 76526 69074 76578
rect 73054 76526 73106 76578
rect 77646 76526 77698 76578
rect 5070 76414 5122 76466
rect 13134 76414 13186 76466
rect 15150 76414 15202 76466
rect 16942 76414 16994 76466
rect 19182 76414 19234 76466
rect 20974 76414 21026 76466
rect 23214 76414 23266 76466
rect 25006 76414 25058 76466
rect 27246 76414 27298 76466
rect 28254 76414 28306 76466
rect 30046 76414 30098 76466
rect 32174 76414 32226 76466
rect 34078 76414 34130 76466
rect 36094 76414 36146 76466
rect 38110 76414 38162 76466
rect 44830 76414 44882 76466
rect 50094 76414 50146 76466
rect 50318 76414 50370 76466
rect 54238 76414 54290 76466
rect 59166 76414 59218 76466
rect 62414 76414 62466 76466
rect 3278 76302 3330 76354
rect 28814 76302 28866 76354
rect 30718 76302 30770 76354
rect 32734 76302 32786 76354
rect 34750 76302 34802 76354
rect 36766 76302 36818 76354
rect 40014 76302 40066 76354
rect 41694 76302 41746 76354
rect 46398 76302 46450 76354
rect 51102 76302 51154 76354
rect 56142 76302 56194 76354
rect 56926 76302 56978 76354
rect 43710 76190 43762 76242
rect 44046 76190 44098 76242
rect 46734 76190 46786 76242
rect 49758 76190 49810 76242
rect 62862 76190 62914 76242
rect 65886 76190 65938 76242
rect 74510 76190 74562 76242
rect 4478 76022 4530 76074
rect 4582 76022 4634 76074
rect 4686 76022 4738 76074
rect 35198 76022 35250 76074
rect 35302 76022 35354 76074
rect 35406 76022 35458 76074
rect 65918 76022 65970 76074
rect 66022 76022 66074 76074
rect 66126 76022 66178 76074
rect 29486 75854 29538 75906
rect 44718 75854 44770 75906
rect 53118 75854 53170 75906
rect 1822 75742 1874 75794
rect 19854 75742 19906 75794
rect 20974 75742 21026 75794
rect 23998 75742 24050 75794
rect 26798 75742 26850 75794
rect 29374 75742 29426 75794
rect 35086 75742 35138 75794
rect 36318 75742 36370 75794
rect 38782 75742 38834 75794
rect 40462 75742 40514 75794
rect 44830 75742 44882 75794
rect 48414 75742 48466 75794
rect 48974 75742 49026 75794
rect 65214 75742 65266 75794
rect 75070 75742 75122 75794
rect 13806 75630 13858 75682
rect 15822 75630 15874 75682
rect 17838 75630 17890 75682
rect 30046 75630 30098 75682
rect 30382 75630 30434 75682
rect 30606 75630 30658 75682
rect 31166 75630 31218 75682
rect 31390 75630 31442 75682
rect 31726 75630 31778 75682
rect 38110 75630 38162 75682
rect 40686 75630 40738 75682
rect 41134 75630 41186 75682
rect 46734 75630 46786 75682
rect 49086 75630 49138 75682
rect 50430 75630 50482 75682
rect 52334 75630 52386 75682
rect 53006 75630 53058 75682
rect 54126 75630 54178 75682
rect 54462 75630 54514 75682
rect 55134 75630 55186 75682
rect 55582 75630 55634 75682
rect 59614 75630 59666 75682
rect 3166 75518 3218 75570
rect 5182 75518 5234 75570
rect 13246 75518 13298 75570
rect 15262 75518 15314 75570
rect 17278 75518 17330 75570
rect 19294 75518 19346 75570
rect 21758 75518 21810 75570
rect 23326 75518 23378 75570
rect 25342 75518 25394 75570
rect 27358 75518 27410 75570
rect 28254 75518 28306 75570
rect 28590 75518 28642 75570
rect 29262 75518 29314 75570
rect 32286 75518 32338 75570
rect 32622 75518 32674 75570
rect 33182 75518 33234 75570
rect 33518 75518 33570 75570
rect 33742 75518 33794 75570
rect 34414 75518 34466 75570
rect 34974 75518 35026 75570
rect 35310 75518 35362 75570
rect 35534 75518 35586 75570
rect 36654 75518 36706 75570
rect 36878 75518 36930 75570
rect 40014 75518 40066 75570
rect 41694 75518 41746 75570
rect 42254 75518 42306 75570
rect 42926 75518 42978 75570
rect 43038 75518 43090 75570
rect 43486 75518 43538 75570
rect 43822 75518 43874 75570
rect 45950 75518 46002 75570
rect 47406 75518 47458 75570
rect 49422 75518 49474 75570
rect 53790 75518 53842 75570
rect 56478 75518 56530 75570
rect 57374 75518 57426 75570
rect 59166 75518 59218 75570
rect 59950 75518 60002 75570
rect 60510 75518 60562 75570
rect 63086 75518 63138 75570
rect 63758 75518 63810 75570
rect 64430 75518 64482 75570
rect 65662 75518 65714 75570
rect 66334 75518 66386 75570
rect 69022 75518 69074 75570
rect 70702 75518 70754 75570
rect 71710 75518 71762 75570
rect 72382 75518 72434 75570
rect 73390 75518 73442 75570
rect 73950 75518 74002 75570
rect 76974 75518 77026 75570
rect 77982 75518 78034 75570
rect 33294 75406 33346 75458
rect 36318 75406 36370 75458
rect 36430 75406 36482 75458
rect 37550 75406 37602 75458
rect 40126 75406 40178 75458
rect 40238 75406 40290 75458
rect 41246 75406 41298 75458
rect 41470 75406 41522 75458
rect 42478 75406 42530 75458
rect 42702 75406 42754 75458
rect 43710 75406 43762 75458
rect 43934 75406 43986 75458
rect 44046 75406 44098 75458
rect 44942 75406 44994 75458
rect 45614 75406 45666 75458
rect 46510 75406 46562 75458
rect 47742 75406 47794 75458
rect 48302 75406 48354 75458
rect 49534 75406 49586 75458
rect 49758 75406 49810 75458
rect 50878 75406 50930 75458
rect 50990 75406 51042 75458
rect 51102 75406 51154 75458
rect 51662 75406 51714 75458
rect 51774 75406 51826 75458
rect 51886 75406 51938 75458
rect 52894 75406 52946 75458
rect 53902 75406 53954 75458
rect 54014 75406 54066 75458
rect 55022 75406 55074 75458
rect 55246 75406 55298 75458
rect 56142 75406 56194 75458
rect 57038 75406 57090 75458
rect 57934 75406 57986 75458
rect 58270 75406 58322 75458
rect 58830 75406 58882 75458
rect 59838 75406 59890 75458
rect 61742 75406 61794 75458
rect 62414 75406 62466 75458
rect 66894 75406 66946 75458
rect 70030 75406 70082 75458
rect 73054 75406 73106 75458
rect 19838 75238 19890 75290
rect 19942 75238 19994 75290
rect 20046 75238 20098 75290
rect 50558 75238 50610 75290
rect 50662 75238 50714 75290
rect 50766 75238 50818 75290
rect 28702 75070 28754 75122
rect 29374 75070 29426 75122
rect 30270 75070 30322 75122
rect 31278 75070 31330 75122
rect 33182 75070 33234 75122
rect 34638 75070 34690 75122
rect 35646 75070 35698 75122
rect 35758 75070 35810 75122
rect 36430 75070 36482 75122
rect 38782 75070 38834 75122
rect 40014 75070 40066 75122
rect 40126 75070 40178 75122
rect 41022 75070 41074 75122
rect 43150 75070 43202 75122
rect 44942 75070 44994 75122
rect 45950 75070 46002 75122
rect 47070 75070 47122 75122
rect 54350 75070 54402 75122
rect 54798 75070 54850 75122
rect 56590 75070 56642 75122
rect 59278 75070 59330 75122
rect 62190 75070 62242 75122
rect 62862 75070 62914 75122
rect 63870 75070 63922 75122
rect 66782 75070 66834 75122
rect 67678 75070 67730 75122
rect 70814 75070 70866 75122
rect 72830 75070 72882 75122
rect 74398 75070 74450 75122
rect 75742 75070 75794 75122
rect 76414 75070 76466 75122
rect 77422 75070 77474 75122
rect 78094 75070 78146 75122
rect 29934 74958 29986 75010
rect 30830 74958 30882 75010
rect 37326 74958 37378 75010
rect 38670 74958 38722 75010
rect 39006 74958 39058 75010
rect 43710 74958 43762 75010
rect 47182 74958 47234 75010
rect 48862 74958 48914 75010
rect 49086 74958 49138 75010
rect 49982 74958 50034 75010
rect 52670 74958 52722 75010
rect 53006 74958 53058 75010
rect 53566 74958 53618 75010
rect 57486 74958 57538 75010
rect 60174 74958 60226 75010
rect 61630 74958 61682 75010
rect 31054 74846 31106 74898
rect 31390 74846 31442 74898
rect 32062 74846 32114 74898
rect 33742 74846 33794 74898
rect 34414 74846 34466 74898
rect 35198 74846 35250 74898
rect 35534 74846 35586 74898
rect 37550 74846 37602 74898
rect 38222 74846 38274 74898
rect 39454 74846 39506 74898
rect 39902 74846 39954 74898
rect 40798 74846 40850 74898
rect 42478 74846 42530 74898
rect 42590 74846 42642 74898
rect 42702 74846 42754 74898
rect 43934 74846 43986 74898
rect 44158 74846 44210 74898
rect 44494 74846 44546 74898
rect 45726 74846 45778 74898
rect 46846 74846 46898 74898
rect 50318 74846 50370 74898
rect 51438 74846 51490 74898
rect 53790 74846 53842 74898
rect 54014 74846 54066 74898
rect 54350 74846 54402 74898
rect 57710 74846 57762 74898
rect 58830 74846 58882 74898
rect 59166 74846 59218 74898
rect 59502 74846 59554 74898
rect 61518 74846 61570 74898
rect 29262 74734 29314 74786
rect 32286 74734 32338 74786
rect 38670 74734 38722 74786
rect 41694 74734 41746 74786
rect 43822 74734 43874 74786
rect 45838 74734 45890 74786
rect 46174 74734 46226 74786
rect 50990 74734 51042 74786
rect 51886 74734 51938 74786
rect 55694 74734 55746 74786
rect 58270 74734 58322 74786
rect 59390 74734 59442 74786
rect 60286 74734 60338 74786
rect 60958 74734 61010 74786
rect 63422 74734 63474 74786
rect 32622 74622 32674 74674
rect 33518 74622 33570 74674
rect 36766 74622 36818 74674
rect 44606 74622 44658 74674
rect 44942 74622 44994 74674
rect 46398 74622 46450 74674
rect 48190 74622 48242 74674
rect 48526 74622 48578 74674
rect 55246 74622 55298 74674
rect 55470 74622 55522 74674
rect 56926 74622 56978 74674
rect 60846 74622 60898 74674
rect 4478 74454 4530 74506
rect 4582 74454 4634 74506
rect 4686 74454 4738 74506
rect 35198 74454 35250 74506
rect 35302 74454 35354 74506
rect 35406 74454 35458 74506
rect 65918 74454 65970 74506
rect 66022 74454 66074 74506
rect 66126 74454 66178 74506
rect 33966 74286 34018 74338
rect 34302 74286 34354 74338
rect 35086 74286 35138 74338
rect 35422 74286 35474 74338
rect 36318 74286 36370 74338
rect 38222 74286 38274 74338
rect 44270 74286 44322 74338
rect 48638 74286 48690 74338
rect 49310 74286 49362 74338
rect 50766 74286 50818 74338
rect 28926 74174 28978 74226
rect 29262 74174 29314 74226
rect 29822 74174 29874 74226
rect 34526 74174 34578 74226
rect 35646 74174 35698 74226
rect 40462 74174 40514 74226
rect 42030 74174 42082 74226
rect 43934 74174 43986 74226
rect 44830 74174 44882 74226
rect 47854 74174 47906 74226
rect 53230 74174 53282 74226
rect 61630 74174 61682 74226
rect 62526 74174 62578 74226
rect 62974 74174 63026 74226
rect 63534 74174 63586 74226
rect 78094 74174 78146 74226
rect 30494 74062 30546 74114
rect 31166 74062 31218 74114
rect 32062 74062 32114 74114
rect 33070 74062 33122 74114
rect 36654 74062 36706 74114
rect 37438 74062 37490 74114
rect 38110 74062 38162 74114
rect 38782 74062 38834 74114
rect 39342 74062 39394 74114
rect 40350 74062 40402 74114
rect 41694 74062 41746 74114
rect 42926 74062 42978 74114
rect 43150 74062 43202 74114
rect 44158 74062 44210 74114
rect 45502 74062 45554 74114
rect 46062 74062 46114 74114
rect 48750 74062 48802 74114
rect 50094 74062 50146 74114
rect 50654 74062 50706 74114
rect 51326 74062 51378 74114
rect 52110 74062 52162 74114
rect 52894 74062 52946 74114
rect 53902 74062 53954 74114
rect 54238 74062 54290 74114
rect 54686 74062 54738 74114
rect 55022 74062 55074 74114
rect 55694 74062 55746 74114
rect 57598 74062 57650 74114
rect 58718 74062 58770 74114
rect 58942 74062 58994 74114
rect 59278 74062 59330 74114
rect 62078 74062 62130 74114
rect 32398 73950 32450 74002
rect 37214 73950 37266 74002
rect 39902 73950 39954 74002
rect 40574 73950 40626 74002
rect 40798 73950 40850 74002
rect 42142 73950 42194 74002
rect 45614 73950 45666 74002
rect 45726 73950 45778 74002
rect 49758 73950 49810 74002
rect 49870 73950 49922 74002
rect 50878 73950 50930 74002
rect 51102 73950 51154 74002
rect 51998 73950 52050 74002
rect 52782 73950 52834 74002
rect 56030 73950 56082 74002
rect 56814 73950 56866 74002
rect 57038 73950 57090 74002
rect 57934 73950 57986 74002
rect 30270 73838 30322 73890
rect 31502 73838 31554 73890
rect 33406 73838 33458 73890
rect 38894 73838 38946 73890
rect 39006 73838 39058 73890
rect 44270 73838 44322 73890
rect 46622 73838 46674 73890
rect 47294 73838 47346 73890
rect 48638 73838 48690 73890
rect 51774 73838 51826 73890
rect 54910 73838 54962 73890
rect 55806 73838 55858 73890
rect 56926 73838 56978 73890
rect 57822 73838 57874 73890
rect 58830 73838 58882 73890
rect 59838 73838 59890 73890
rect 60510 73838 60562 73890
rect 19838 73670 19890 73722
rect 19942 73670 19994 73722
rect 20046 73670 20098 73722
rect 50558 73670 50610 73722
rect 50662 73670 50714 73722
rect 50766 73670 50818 73722
rect 30942 73502 30994 73554
rect 31390 73502 31442 73554
rect 32174 73502 32226 73554
rect 32734 73502 32786 73554
rect 33406 73502 33458 73554
rect 33518 73502 33570 73554
rect 34526 73502 34578 73554
rect 35422 73502 35474 73554
rect 36318 73502 36370 73554
rect 36654 73502 36706 73554
rect 36878 73502 36930 73554
rect 39678 73502 39730 73554
rect 40910 73502 40962 73554
rect 42254 73502 42306 73554
rect 47854 73502 47906 73554
rect 48526 73502 48578 73554
rect 50318 73502 50370 73554
rect 54574 73502 54626 73554
rect 55358 73502 55410 73554
rect 55918 73502 55970 73554
rect 56030 73502 56082 73554
rect 60398 73502 60450 73554
rect 60958 73502 61010 73554
rect 61406 73502 61458 73554
rect 61854 73502 61906 73554
rect 33630 73390 33682 73442
rect 34190 73390 34242 73442
rect 35310 73390 35362 73442
rect 35982 73390 36034 73442
rect 36094 73390 36146 73442
rect 37550 73390 37602 73442
rect 37886 73390 37938 73442
rect 40574 73390 40626 73442
rect 44606 73390 44658 73442
rect 44718 73390 44770 73442
rect 47182 73390 47234 73442
rect 50878 73390 50930 73442
rect 51102 73390 51154 73442
rect 52894 73390 52946 73442
rect 54014 73390 54066 73442
rect 54910 73390 54962 73442
rect 57262 73390 57314 73442
rect 36990 73278 37042 73330
rect 38446 73278 38498 73330
rect 40798 73278 40850 73330
rect 41022 73278 41074 73330
rect 43150 73278 43202 73330
rect 44158 73278 44210 73330
rect 44382 73278 44434 73330
rect 45950 73278 46002 73330
rect 47294 73278 47346 73330
rect 51214 73278 51266 73330
rect 51550 73278 51602 73330
rect 52446 73278 52498 73330
rect 53566 73278 53618 73330
rect 53678 73278 53730 73330
rect 53902 73278 53954 73330
rect 56142 73278 56194 73330
rect 56590 73278 56642 73330
rect 57710 73278 57762 73330
rect 59278 73278 59330 73330
rect 30382 73166 30434 73218
rect 39790 73166 39842 73218
rect 41694 73166 41746 73218
rect 42702 73166 42754 73218
rect 45502 73166 45554 73218
rect 45838 73166 45890 73218
rect 47966 73166 48018 73218
rect 49422 73166 49474 73218
rect 50766 73166 50818 73218
rect 52110 73166 52162 73218
rect 58046 73166 58098 73218
rect 58830 73166 58882 73218
rect 59614 73166 59666 73218
rect 38670 73054 38722 73106
rect 39006 73054 39058 73106
rect 39902 73054 39954 73106
rect 42926 73054 42978 73106
rect 44942 73054 44994 73106
rect 47182 73054 47234 73106
rect 49646 73054 49698 73106
rect 49870 73054 49922 73106
rect 4478 72886 4530 72938
rect 4582 72886 4634 72938
rect 4686 72886 4738 72938
rect 35198 72886 35250 72938
rect 35302 72886 35354 72938
rect 35406 72886 35458 72938
rect 65918 72886 65970 72938
rect 66022 72886 66074 72938
rect 66126 72886 66178 72938
rect 33742 72718 33794 72770
rect 34302 72718 34354 72770
rect 55582 72718 55634 72770
rect 57150 72718 57202 72770
rect 31950 72606 32002 72658
rect 32398 72606 32450 72658
rect 32846 72606 32898 72658
rect 33294 72606 33346 72658
rect 33742 72606 33794 72658
rect 34190 72606 34242 72658
rect 35422 72606 35474 72658
rect 36990 72606 37042 72658
rect 43150 72606 43202 72658
rect 43934 72606 43986 72658
rect 45614 72606 45666 72658
rect 49758 72606 49810 72658
rect 50878 72606 50930 72658
rect 51550 72606 51602 72658
rect 54910 72606 54962 72658
rect 56478 72606 56530 72658
rect 58046 72606 58098 72658
rect 59278 72606 59330 72658
rect 59726 72606 59778 72658
rect 60174 72606 60226 72658
rect 60622 72606 60674 72658
rect 37438 72494 37490 72546
rect 37886 72494 37938 72546
rect 39006 72494 39058 72546
rect 39678 72494 39730 72546
rect 39902 72494 39954 72546
rect 40350 72494 40402 72546
rect 40574 72494 40626 72546
rect 42814 72494 42866 72546
rect 45166 72494 45218 72546
rect 46286 72494 46338 72546
rect 46622 72494 46674 72546
rect 49646 72494 49698 72546
rect 49870 72494 49922 72546
rect 50766 72494 50818 72546
rect 51886 72494 51938 72546
rect 52446 72494 52498 72546
rect 53342 72494 53394 72546
rect 54686 72494 54738 72546
rect 55694 72494 55746 72546
rect 57038 72494 57090 72546
rect 57262 72494 57314 72546
rect 57934 72494 57986 72546
rect 34750 72382 34802 72434
rect 36430 72382 36482 72434
rect 40238 72382 40290 72434
rect 42254 72382 42306 72434
rect 43934 72382 43986 72434
rect 44158 72382 44210 72434
rect 44718 72382 44770 72434
rect 46398 72382 46450 72434
rect 47070 72382 47122 72434
rect 48190 72382 48242 72434
rect 49086 72382 49138 72434
rect 50094 72382 50146 72434
rect 51662 72382 51714 72434
rect 52670 72382 52722 72434
rect 54350 72382 54402 72434
rect 55582 72382 55634 72434
rect 59166 72382 59218 72434
rect 35310 72270 35362 72322
rect 38558 72270 38610 72322
rect 41694 72270 41746 72322
rect 47630 72270 47682 72322
rect 19838 72102 19890 72154
rect 19942 72102 19994 72154
rect 20046 72102 20098 72154
rect 50558 72102 50610 72154
rect 50662 72102 50714 72154
rect 50766 72102 50818 72154
rect 33854 71934 33906 71986
rect 35982 71934 36034 71986
rect 36430 71934 36482 71986
rect 36990 71934 37042 71986
rect 37438 71934 37490 71986
rect 37662 71934 37714 71986
rect 38446 71934 38498 71986
rect 41022 71934 41074 71986
rect 43038 71934 43090 71986
rect 45726 71934 45778 71986
rect 47182 71934 47234 71986
rect 47630 71934 47682 71986
rect 48078 71934 48130 71986
rect 52334 71934 52386 71986
rect 54462 71934 54514 71986
rect 58046 71934 58098 71986
rect 58718 71934 58770 71986
rect 59278 71934 59330 71986
rect 59614 71934 59666 71986
rect 37774 71822 37826 71874
rect 40126 71822 40178 71874
rect 43262 71822 43314 71874
rect 43934 71822 43986 71874
rect 45166 71822 45218 71874
rect 49422 71822 49474 71874
rect 53006 71822 53058 71874
rect 55470 71822 55522 71874
rect 56702 71822 56754 71874
rect 57934 71822 57986 71874
rect 39006 71710 39058 71762
rect 39790 71710 39842 71762
rect 41806 71710 41858 71762
rect 42814 71710 42866 71762
rect 43598 71710 43650 71762
rect 44494 71710 44546 71762
rect 44942 71710 44994 71762
rect 45950 71710 46002 71762
rect 46174 71710 46226 71762
rect 50206 71710 50258 71762
rect 51550 71710 51602 71762
rect 53230 71710 53282 71762
rect 53566 71710 53618 71762
rect 55246 71710 55298 71762
rect 56926 71710 56978 71762
rect 34974 71598 35026 71650
rect 35422 71598 35474 71650
rect 44718 71598 44770 71650
rect 46286 71598 46338 71650
rect 46734 71598 46786 71650
rect 48526 71598 48578 71650
rect 51662 71598 51714 71650
rect 34862 71486 34914 71538
rect 46062 71486 46114 71538
rect 46734 71486 46786 71538
rect 47966 71486 48018 71538
rect 48526 71486 48578 71538
rect 4478 71318 4530 71370
rect 4582 71318 4634 71370
rect 4686 71318 4738 71370
rect 35198 71318 35250 71370
rect 35302 71318 35354 71370
rect 35406 71318 35458 71370
rect 65918 71318 65970 71370
rect 66022 71318 66074 71370
rect 66126 71318 66178 71370
rect 39902 71150 39954 71202
rect 41582 71150 41634 71202
rect 45614 71150 45666 71202
rect 46286 71150 46338 71202
rect 46510 71150 46562 71202
rect 46958 71150 47010 71202
rect 54462 71150 54514 71202
rect 54686 71150 54738 71202
rect 54910 71150 54962 71202
rect 56142 71150 56194 71202
rect 56478 71150 56530 71202
rect 57374 71150 57426 71202
rect 35198 71038 35250 71090
rect 35646 71038 35698 71090
rect 37326 71038 37378 71090
rect 37662 71038 37714 71090
rect 38222 71038 38274 71090
rect 40910 71038 40962 71090
rect 42142 71038 42194 71090
rect 45614 71038 45666 71090
rect 46062 71038 46114 71090
rect 46958 71038 47010 71090
rect 47406 71038 47458 71090
rect 47854 71038 47906 71090
rect 48750 71038 48802 71090
rect 49310 71038 49362 71090
rect 50878 71038 50930 71090
rect 51326 71038 51378 71090
rect 51886 71038 51938 71090
rect 52894 71038 52946 71090
rect 53230 71038 53282 71090
rect 54126 71038 54178 71090
rect 54462 71038 54514 71090
rect 54910 71038 54962 71090
rect 57262 71038 57314 71090
rect 57934 71038 57986 71090
rect 36430 70926 36482 70978
rect 39006 70926 39058 70978
rect 41134 70926 41186 70978
rect 42814 70926 42866 70978
rect 43598 70926 43650 70978
rect 44270 70926 44322 70978
rect 44942 70926 44994 70978
rect 46510 70926 46562 70978
rect 51774 70926 51826 70978
rect 52110 70926 52162 70978
rect 52334 70926 52386 70978
rect 55918 70926 55970 70978
rect 57038 70926 57090 70978
rect 38670 70814 38722 70866
rect 39790 70814 39842 70866
rect 50206 70814 50258 70866
rect 36094 70702 36146 70754
rect 39902 70702 39954 70754
rect 48302 70702 48354 70754
rect 49646 70702 49698 70754
rect 55470 70702 55522 70754
rect 19838 70534 19890 70586
rect 19942 70534 19994 70586
rect 20046 70534 20098 70586
rect 50558 70534 50610 70586
rect 50662 70534 50714 70586
rect 50766 70534 50818 70586
rect 38110 70366 38162 70418
rect 38558 70366 38610 70418
rect 39006 70366 39058 70418
rect 39454 70366 39506 70418
rect 40126 70366 40178 70418
rect 40350 70366 40402 70418
rect 41022 70366 41074 70418
rect 42814 70366 42866 70418
rect 43934 70366 43986 70418
rect 44270 70366 44322 70418
rect 44830 70366 44882 70418
rect 45278 70366 45330 70418
rect 45726 70366 45778 70418
rect 46174 70366 46226 70418
rect 46622 70366 46674 70418
rect 47182 70366 47234 70418
rect 49758 70366 49810 70418
rect 50206 70366 50258 70418
rect 50654 70366 50706 70418
rect 51102 70366 51154 70418
rect 51662 70366 51714 70418
rect 52558 70366 52610 70418
rect 53006 70366 53058 70418
rect 54238 70366 54290 70418
rect 54686 70366 54738 70418
rect 55358 70366 55410 70418
rect 56030 70366 56082 70418
rect 56478 70366 56530 70418
rect 40462 70254 40514 70306
rect 56926 70254 56978 70306
rect 37214 70142 37266 70194
rect 37550 70142 37602 70194
rect 43150 70142 43202 70194
rect 43374 70142 43426 70194
rect 39566 70030 39618 70082
rect 53454 70030 53506 70082
rect 37998 69918 38050 69970
rect 38558 69918 38610 69970
rect 43710 69918 43762 69970
rect 44718 69918 44770 69970
rect 4478 69750 4530 69802
rect 4582 69750 4634 69802
rect 4686 69750 4738 69802
rect 35198 69750 35250 69802
rect 35302 69750 35354 69802
rect 35406 69750 35458 69802
rect 65918 69750 65970 69802
rect 66022 69750 66074 69802
rect 66126 69750 66178 69802
rect 38558 69470 38610 69522
rect 39006 69470 39058 69522
rect 39678 69470 39730 69522
rect 40126 69470 40178 69522
rect 43262 69470 43314 69522
rect 44494 69470 44546 69522
rect 44830 69470 44882 69522
rect 54686 69470 54738 69522
rect 19838 68966 19890 69018
rect 19942 68966 19994 69018
rect 20046 68966 20098 69018
rect 50558 68966 50610 69018
rect 50662 68966 50714 69018
rect 50766 68966 50818 69018
rect 4478 68182 4530 68234
rect 4582 68182 4634 68234
rect 4686 68182 4738 68234
rect 35198 68182 35250 68234
rect 35302 68182 35354 68234
rect 35406 68182 35458 68234
rect 65918 68182 65970 68234
rect 66022 68182 66074 68234
rect 66126 68182 66178 68234
rect 19838 67398 19890 67450
rect 19942 67398 19994 67450
rect 20046 67398 20098 67450
rect 50558 67398 50610 67450
rect 50662 67398 50714 67450
rect 50766 67398 50818 67450
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 35198 66614 35250 66666
rect 35302 66614 35354 66666
rect 35406 66614 35458 66666
rect 65918 66614 65970 66666
rect 66022 66614 66074 66666
rect 66126 66614 66178 66666
rect 19838 65830 19890 65882
rect 19942 65830 19994 65882
rect 20046 65830 20098 65882
rect 50558 65830 50610 65882
rect 50662 65830 50714 65882
rect 50766 65830 50818 65882
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 35198 65046 35250 65098
rect 35302 65046 35354 65098
rect 35406 65046 35458 65098
rect 65918 65046 65970 65098
rect 66022 65046 66074 65098
rect 66126 65046 66178 65098
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 50558 64262 50610 64314
rect 50662 64262 50714 64314
rect 50766 64262 50818 64314
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 65918 63478 65970 63530
rect 66022 63478 66074 63530
rect 66126 63478 66178 63530
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 50558 62694 50610 62746
rect 50662 62694 50714 62746
rect 50766 62694 50818 62746
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 65918 61910 65970 61962
rect 66022 61910 66074 61962
rect 66126 61910 66178 61962
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 50558 61126 50610 61178
rect 50662 61126 50714 61178
rect 50766 61126 50818 61178
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 65918 60342 65970 60394
rect 66022 60342 66074 60394
rect 66126 60342 66178 60394
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 50558 59558 50610 59610
rect 50662 59558 50714 59610
rect 50766 59558 50818 59610
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 65918 58774 65970 58826
rect 66022 58774 66074 58826
rect 66126 58774 66178 58826
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 50558 57990 50610 58042
rect 50662 57990 50714 58042
rect 50766 57990 50818 58042
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 65918 57206 65970 57258
rect 66022 57206 66074 57258
rect 66126 57206 66178 57258
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 65918 55638 65970 55690
rect 66022 55638 66074 55690
rect 66126 55638 66178 55690
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 65918 54070 65970 54122
rect 66022 54070 66074 54122
rect 66126 54070 66178 54122
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 65918 52502 65970 52554
rect 66022 52502 66074 52554
rect 66126 52502 66178 52554
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 65918 50934 65970 50986
rect 66022 50934 66074 50986
rect 66126 50934 66178 50986
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 65918 49366 65970 49418
rect 66022 49366 66074 49418
rect 66126 49366 66178 49418
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 65918 47798 65970 47850
rect 66022 47798 66074 47850
rect 66126 47798 66178 47850
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 65918 46230 65970 46282
rect 66022 46230 66074 46282
rect 66126 46230 66178 46282
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 65918 44662 65970 44714
rect 66022 44662 66074 44714
rect 66126 44662 66178 44714
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 65918 43094 65970 43146
rect 66022 43094 66074 43146
rect 66126 43094 66178 43146
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 65918 41526 65970 41578
rect 66022 41526 66074 41578
rect 66126 41526 66178 41578
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 65918 39958 65970 40010
rect 66022 39958 66074 40010
rect 66126 39958 66178 40010
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 65918 38390 65970 38442
rect 66022 38390 66074 38442
rect 66126 38390 66178 38442
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 65918 36822 65970 36874
rect 66022 36822 66074 36874
rect 66126 36822 66178 36874
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 65918 35254 65970 35306
rect 66022 35254 66074 35306
rect 66126 35254 66178 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 65918 33686 65970 33738
rect 66022 33686 66074 33738
rect 66126 33686 66178 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 65918 32118 65970 32170
rect 66022 32118 66074 32170
rect 66126 32118 66178 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 65918 30550 65970 30602
rect 66022 30550 66074 30602
rect 66126 30550 66178 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 65918 28982 65970 29034
rect 66022 28982 66074 29034
rect 66126 28982 66178 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 65918 27414 65970 27466
rect 66022 27414 66074 27466
rect 66126 27414 66178 27466
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 65918 25846 65970 25898
rect 66022 25846 66074 25898
rect 66126 25846 66178 25898
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 65918 24278 65970 24330
rect 66022 24278 66074 24330
rect 66126 24278 66178 24330
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 65918 22710 65970 22762
rect 66022 22710 66074 22762
rect 66126 22710 66178 22762
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 65918 21142 65970 21194
rect 66022 21142 66074 21194
rect 66126 21142 66178 21194
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 65918 19574 65970 19626
rect 66022 19574 66074 19626
rect 66126 19574 66178 19626
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 65918 18006 65970 18058
rect 66022 18006 66074 18058
rect 66126 18006 66178 18058
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 65918 16438 65970 16490
rect 66022 16438 66074 16490
rect 66126 16438 66178 16490
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 65918 14870 65970 14922
rect 66022 14870 66074 14922
rect 66126 14870 66178 14922
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 65918 13302 65970 13354
rect 66022 13302 66074 13354
rect 66126 13302 66178 13354
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 65918 11734 65970 11786
rect 66022 11734 66074 11786
rect 66126 11734 66178 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 65918 10166 65970 10218
rect 66022 10166 66074 10218
rect 66126 10166 66178 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 65918 8598 65970 8650
rect 66022 8598 66074 8650
rect 66126 8598 66178 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 65918 7030 65970 7082
rect 66022 7030 66074 7082
rect 66126 7030 66178 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 65918 5462 65970 5514
rect 66022 5462 66074 5514
rect 66126 5462 66178 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 73278 4398 73330 4450
rect 73950 4398 74002 4450
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 65918 3894 65970 3946
rect 66022 3894 66074 3946
rect 66126 3894 66178 3946
rect 6974 3278 7026 3330
rect 8318 3278 8370 3330
rect 9214 3278 9266 3330
rect 10110 3278 10162 3330
rect 10782 3278 10834 3330
rect 11566 3278 11618 3330
rect 12238 3278 12290 3330
rect 12910 3278 12962 3330
rect 13582 3278 13634 3330
rect 14254 3278 14306 3330
rect 14926 3278 14978 3330
rect 15598 3278 15650 3330
rect 16270 3278 16322 3330
rect 16942 3278 16994 3330
rect 17614 3278 17666 3330
rect 18286 3278 18338 3330
rect 18958 3278 19010 3330
rect 19630 3278 19682 3330
rect 20302 3278 20354 3330
rect 20974 3278 21026 3330
rect 21758 3278 21810 3330
rect 22430 3278 22482 3330
rect 23102 3278 23154 3330
rect 23774 3278 23826 3330
rect 24446 3278 24498 3330
rect 25118 3278 25170 3330
rect 25790 3278 25842 3330
rect 26462 3278 26514 3330
rect 27134 3278 27186 3330
rect 27806 3278 27858 3330
rect 28478 3278 28530 3330
rect 29150 3278 29202 3330
rect 29822 3278 29874 3330
rect 30494 3278 30546 3330
rect 31166 3278 31218 3330
rect 31838 3278 31890 3330
rect 32510 3278 32562 3330
rect 33182 3278 33234 3330
rect 33854 3278 33906 3330
rect 34526 3278 34578 3330
rect 35198 3278 35250 3330
rect 35870 3278 35922 3330
rect 36542 3278 36594 3330
rect 37214 3278 37266 3330
rect 37886 3278 37938 3330
rect 38558 3278 38610 3330
rect 39230 3278 39282 3330
rect 39902 3278 39954 3330
rect 40574 3278 40626 3330
rect 41694 3278 41746 3330
rect 42366 3278 42418 3330
rect 43038 3278 43090 3330
rect 43710 3278 43762 3330
rect 44382 3278 44434 3330
rect 45054 3278 45106 3330
rect 45726 3278 45778 3330
rect 46398 3278 46450 3330
rect 47070 3278 47122 3330
rect 47742 3278 47794 3330
rect 48414 3278 48466 3330
rect 49086 3278 49138 3330
rect 49758 3278 49810 3330
rect 50430 3278 50482 3330
rect 51102 3278 51154 3330
rect 51774 3278 51826 3330
rect 52446 3278 52498 3330
rect 53118 3278 53170 3330
rect 53790 3278 53842 3330
rect 54462 3278 54514 3330
rect 55134 3278 55186 3330
rect 55806 3278 55858 3330
rect 56478 3278 56530 3330
rect 57150 3278 57202 3330
rect 57822 3278 57874 3330
rect 58494 3278 58546 3330
rect 59166 3278 59218 3330
rect 59838 3278 59890 3330
rect 60510 3278 60562 3330
rect 61630 3278 61682 3330
rect 62302 3278 62354 3330
rect 62974 3278 63026 3330
rect 63646 3278 63698 3330
rect 64318 3278 64370 3330
rect 64990 3278 65042 3330
rect 65662 3278 65714 3330
rect 66334 3278 66386 3330
rect 67006 3278 67058 3330
rect 67678 3278 67730 3330
rect 68350 3278 68402 3330
rect 69022 3278 69074 3330
rect 69694 3278 69746 3330
rect 70366 3278 70418 3330
rect 71038 3278 71090 3330
rect 71710 3278 71762 3330
rect 72382 3278 72434 3330
rect 73054 3278 73106 3330
rect 73726 3278 73778 3330
rect 74398 3278 74450 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
rect 54574 1934 54626 1986
rect 55134 1934 55186 1986
rect 42366 1822 42418 1874
rect 43038 1822 43090 1874
rect 44494 1822 44546 1874
rect 45054 1822 45106 1874
rect 47854 1822 47906 1874
rect 48414 1822 48466 1874
rect 51214 1822 51266 1874
rect 51774 1822 51826 1874
rect 57934 1822 57986 1874
rect 58494 1822 58546 1874
rect 41022 1710 41074 1762
rect 41694 1710 41746 1762
rect 43710 1710 43762 1762
rect 44382 1710 44434 1762
rect 45726 1710 45778 1762
rect 46398 1710 46450 1762
rect 47070 1710 47122 1762
rect 47742 1710 47794 1762
rect 49086 1710 49138 1762
rect 49758 1710 49810 1762
rect 50430 1710 50482 1762
rect 51102 1710 51154 1762
rect 52446 1710 52498 1762
rect 53118 1710 53170 1762
rect 53790 1710 53842 1762
rect 54462 1710 54514 1762
rect 55918 1710 55970 1762
rect 56478 1710 56530 1762
rect 57150 1710 57202 1762
rect 57822 1710 57874 1762
rect 59166 1710 59218 1762
rect 59838 1710 59890 1762
rect 60510 1710 60562 1762
rect 61630 1710 61682 1762
rect 62526 1710 62578 1762
rect 63646 1710 63698 1762
rect 63870 1710 63922 1762
rect 64990 1710 65042 1762
rect 65886 1710 65938 1762
rect 67006 1710 67058 1762
rect 67230 1710 67282 1762
rect 68350 1710 68402 1762
rect 69246 1710 69298 1762
rect 70366 1710 70418 1762
rect 70590 1710 70642 1762
rect 71710 1710 71762 1762
rect 72606 1710 72658 1762
rect 73726 1710 73778 1762
<< metal2 >>
rect 1568 79200 1680 80000
rect 2240 79200 2352 80000
rect 2912 79200 3024 80000
rect 3584 79200 3696 80000
rect 4256 79200 4368 80000
rect 4928 79200 5040 80000
rect 5600 79200 5712 80000
rect 6272 79200 6384 80000
rect 6944 79200 7056 80000
rect 7616 79200 7728 80000
rect 8288 79200 8400 80000
rect 8960 79200 9072 80000
rect 9632 79200 9744 80000
rect 10304 79200 10416 80000
rect 10976 79200 11088 80000
rect 11648 79200 11760 80000
rect 12320 79200 12432 80000
rect 12992 79200 13104 80000
rect 13664 79200 13776 80000
rect 14336 79200 14448 80000
rect 15008 79200 15120 80000
rect 15680 79200 15792 80000
rect 16352 79200 16464 80000
rect 17024 79200 17136 80000
rect 17696 79200 17808 80000
rect 18368 79200 18480 80000
rect 19040 79200 19152 80000
rect 19712 79200 19824 80000
rect 20384 79200 20496 80000
rect 21056 79200 21168 80000
rect 21728 79200 21840 80000
rect 22400 79200 22512 80000
rect 23072 79200 23184 80000
rect 23744 79200 23856 80000
rect 24416 79200 24528 80000
rect 25088 79200 25200 80000
rect 25760 79200 25872 80000
rect 26432 79200 26544 80000
rect 27104 79200 27216 80000
rect 27776 79200 27888 80000
rect 28448 79200 28560 80000
rect 29120 79200 29232 80000
rect 29792 79200 29904 80000
rect 30464 79200 30576 80000
rect 31136 79200 31248 80000
rect 31808 79200 31920 80000
rect 32480 79200 32592 80000
rect 33152 79200 33264 80000
rect 33824 79200 33936 80000
rect 34496 79200 34608 80000
rect 35168 79200 35280 80000
rect 35840 79200 35952 80000
rect 36512 79200 36624 80000
rect 37184 79200 37296 80000
rect 37856 79200 37968 80000
rect 38528 79200 38640 80000
rect 39200 79200 39312 80000
rect 39872 79200 39984 80000
rect 40544 79200 40656 80000
rect 41216 79200 41328 80000
rect 41888 79200 42000 80000
rect 42560 79200 42672 80000
rect 43232 79200 43344 80000
rect 43904 79200 44016 80000
rect 44576 79200 44688 80000
rect 45248 79200 45360 80000
rect 45920 79200 46032 80000
rect 46592 79200 46704 80000
rect 47264 79200 47376 80000
rect 47936 79200 48048 80000
rect 48608 79200 48720 80000
rect 49280 79200 49392 80000
rect 49952 79200 50064 80000
rect 50624 79200 50736 80000
rect 51296 79200 51408 80000
rect 51968 79200 52080 80000
rect 52640 79200 52752 80000
rect 53312 79200 53424 80000
rect 53984 79200 54096 80000
rect 54656 79200 54768 80000
rect 55328 79200 55440 80000
rect 56000 79200 56112 80000
rect 56672 79200 56784 80000
rect 57344 79200 57456 80000
rect 58016 79200 58128 80000
rect 58688 79200 58800 80000
rect 59360 79200 59472 80000
rect 60032 79200 60144 80000
rect 60704 79200 60816 80000
rect 61376 79200 61488 80000
rect 62048 79200 62160 80000
rect 62720 79200 62832 80000
rect 63392 79200 63504 80000
rect 64064 79200 64176 80000
rect 64736 79200 64848 80000
rect 65408 79200 65520 80000
rect 66080 79200 66192 80000
rect 66752 79200 66864 80000
rect 67424 79200 67536 80000
rect 68096 79200 68208 80000
rect 68768 79200 68880 80000
rect 69440 79200 69552 80000
rect 70112 79200 70224 80000
rect 70784 79200 70896 80000
rect 71456 79200 71568 80000
rect 72128 79200 72240 80000
rect 72800 79200 72912 80000
rect 73472 79200 73584 80000
rect 74144 79200 74256 80000
rect 74816 79200 74928 80000
rect 75488 79200 75600 80000
rect 76160 79200 76272 80000
rect 76832 79200 76944 80000
rect 77504 79200 77616 80000
rect 78176 79200 78288 80000
rect 1596 76580 1652 79200
rect 1932 76580 1988 76590
rect 1596 76578 1988 76580
rect 1596 76526 1934 76578
rect 1986 76526 1988 76578
rect 1596 76524 1988 76526
rect 1820 75794 1876 76524
rect 1932 76514 1988 76524
rect 1820 75742 1822 75794
rect 1874 75742 1876 75794
rect 1820 75730 1876 75742
rect 2940 75572 2996 79200
rect 3612 76580 3668 79200
rect 3948 76580 4004 76590
rect 3612 76578 4004 76580
rect 3612 76526 3950 76578
rect 4002 76526 4004 76578
rect 3612 76524 4004 76526
rect 3948 76514 4004 76524
rect 3276 76356 3332 76366
rect 3276 76354 3444 76356
rect 3276 76302 3278 76354
rect 3330 76302 3444 76354
rect 3276 76300 3444 76302
rect 3276 76290 3332 76300
rect 3388 75908 3444 76300
rect 4476 76076 4740 76086
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4476 76010 4740 76020
rect 3388 75842 3444 75852
rect 3164 75572 3220 75582
rect 2940 75570 3220 75572
rect 2940 75518 3166 75570
rect 3218 75518 3220 75570
rect 2940 75516 3220 75518
rect 4956 75572 5012 79200
rect 5628 76692 5684 79200
rect 6524 77364 6580 77374
rect 5852 76692 5908 76702
rect 5628 76690 5908 76692
rect 5628 76638 5854 76690
rect 5906 76638 5908 76690
rect 5628 76636 5908 76638
rect 5852 76626 5908 76636
rect 6524 76690 6580 77308
rect 6524 76638 6526 76690
rect 6578 76638 6580 76690
rect 5068 76468 5124 76478
rect 5068 76374 5124 76412
rect 6524 76468 6580 76638
rect 6972 76692 7028 79200
rect 7196 76692 7252 76702
rect 6972 76690 7252 76692
rect 6972 76638 7198 76690
rect 7250 76638 7252 76690
rect 6972 76636 7252 76638
rect 7644 76692 7700 79200
rect 7868 76692 7924 76702
rect 7644 76690 7924 76692
rect 7644 76638 7870 76690
rect 7922 76638 7924 76690
rect 7644 76636 7924 76638
rect 8988 76692 9044 79200
rect 9212 76692 9268 76702
rect 8988 76690 9268 76692
rect 8988 76638 9214 76690
rect 9266 76638 9268 76690
rect 8988 76636 9268 76638
rect 9660 76692 9716 79200
rect 9884 76692 9940 76702
rect 9660 76690 9940 76692
rect 9660 76638 9886 76690
rect 9938 76638 9940 76690
rect 9660 76636 9940 76638
rect 11004 76692 11060 79200
rect 11228 76692 11284 76702
rect 11004 76690 11284 76692
rect 11004 76638 11230 76690
rect 11282 76638 11284 76690
rect 11004 76636 11284 76638
rect 7196 76626 7252 76636
rect 7868 76626 7924 76636
rect 9212 76626 9268 76636
rect 9884 76626 9940 76636
rect 11228 76626 11284 76636
rect 11676 76580 11732 79200
rect 12012 76580 12068 76590
rect 11676 76578 12068 76580
rect 11676 76526 12014 76578
rect 12066 76526 12068 76578
rect 11676 76524 12068 76526
rect 12012 76514 12068 76524
rect 6524 76402 6580 76412
rect 5180 75572 5236 75582
rect 4956 75570 5236 75572
rect 4956 75518 5182 75570
rect 5234 75518 5236 75570
rect 4956 75516 5236 75518
rect 13020 75572 13076 79200
rect 13692 77812 13748 79200
rect 13692 77756 14084 77812
rect 14028 76578 14084 77756
rect 14028 76526 14030 76578
rect 14082 76526 14084 76578
rect 14028 76514 14084 76526
rect 13132 76468 13188 76478
rect 13132 76374 13188 76412
rect 13804 76468 13860 76478
rect 13804 75682 13860 76412
rect 13804 75630 13806 75682
rect 13858 75630 13860 75682
rect 13244 75572 13300 75582
rect 13020 75570 13300 75572
rect 13020 75518 13246 75570
rect 13298 75518 13300 75570
rect 13020 75516 13300 75518
rect 3164 75506 3220 75516
rect 5180 75506 5236 75516
rect 13244 75506 13300 75516
rect 4476 74508 4740 74518
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4476 74442 4740 74452
rect 4476 72940 4740 72950
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4476 72874 4740 72884
rect 13804 71540 13860 75630
rect 15036 75572 15092 79200
rect 15708 77812 15764 79200
rect 15708 77756 16100 77812
rect 16044 76578 16100 77756
rect 16044 76526 16046 76578
rect 16098 76526 16100 76578
rect 16044 76514 16100 76526
rect 15148 76468 15204 76478
rect 15148 76374 15204 76412
rect 15820 76468 15876 76478
rect 15820 75682 15876 76412
rect 15820 75630 15822 75682
rect 15874 75630 15876 75682
rect 15260 75572 15316 75582
rect 15036 75570 15316 75572
rect 15036 75518 15262 75570
rect 15314 75518 15316 75570
rect 15036 75516 15316 75518
rect 15260 75506 15316 75516
rect 15820 72324 15876 75630
rect 16940 76466 16996 76478
rect 16940 76414 16942 76466
rect 16994 76414 16996 76466
rect 16940 75684 16996 76414
rect 16940 75618 16996 75628
rect 17052 75572 17108 79200
rect 17724 76580 17780 79200
rect 18060 76580 18116 76590
rect 17724 76578 18116 76580
rect 17724 76526 18062 76578
rect 18114 76526 18116 76578
rect 17724 76524 18116 76526
rect 18060 76514 18116 76524
rect 17836 75684 17892 75694
rect 17836 75590 17892 75628
rect 17276 75572 17332 75582
rect 17052 75570 17332 75572
rect 17052 75518 17278 75570
rect 17330 75518 17332 75570
rect 17052 75516 17332 75518
rect 19068 75572 19124 79200
rect 19740 77700 19796 79200
rect 19628 77644 19796 77700
rect 19628 76692 19684 77644
rect 19836 76860 20100 76870
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 19836 76794 20100 76804
rect 19628 76636 19908 76692
rect 19852 76578 19908 76636
rect 19852 76526 19854 76578
rect 19906 76526 19908 76578
rect 19852 76514 19908 76526
rect 19180 76466 19236 76478
rect 19180 76414 19182 76466
rect 19234 76414 19236 76466
rect 19180 75796 19236 76414
rect 20972 76466 21028 76478
rect 20972 76414 20974 76466
rect 21026 76414 21028 76466
rect 20972 76244 21028 76414
rect 19180 75730 19236 75740
rect 19852 75796 19908 75806
rect 19852 75684 19908 75740
rect 20972 75794 21028 76188
rect 20972 75742 20974 75794
rect 21026 75742 21028 75794
rect 20972 75730 21028 75742
rect 19852 75628 20244 75684
rect 19292 75572 19348 75582
rect 19068 75570 19348 75572
rect 19068 75518 19294 75570
rect 19346 75518 19348 75570
rect 19068 75516 19348 75518
rect 17276 75506 17332 75516
rect 19292 75506 19348 75516
rect 19836 75292 20100 75302
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 19836 75226 20100 75236
rect 20188 75124 20244 75628
rect 21084 75572 21140 79200
rect 21756 76580 21812 79200
rect 22092 76580 22148 76590
rect 21756 76578 22148 76580
rect 21756 76526 22094 76578
rect 22146 76526 22148 76578
rect 21756 76524 22148 76526
rect 22092 76514 22148 76524
rect 21084 75506 21140 75516
rect 21644 75908 21700 75918
rect 20188 75058 20244 75068
rect 21644 75012 21700 75852
rect 21756 75572 21812 75582
rect 23100 75572 23156 79200
rect 23772 76580 23828 79200
rect 24108 76580 24164 76590
rect 23772 76578 24164 76580
rect 23772 76526 24110 76578
rect 24162 76526 24164 76578
rect 23772 76524 24164 76526
rect 24108 76514 24164 76524
rect 23212 76466 23268 76478
rect 23212 76414 23214 76466
rect 23266 76414 23268 76466
rect 23212 76132 23268 76414
rect 25004 76468 25060 76478
rect 25004 76374 25060 76412
rect 23212 76066 23268 76076
rect 23996 76132 24052 76142
rect 23996 75794 24052 76076
rect 23996 75742 23998 75794
rect 24050 75742 24052 75794
rect 23996 75730 24052 75742
rect 23324 75572 23380 75582
rect 23100 75570 23380 75572
rect 23100 75518 23326 75570
rect 23378 75518 23380 75570
rect 23100 75516 23380 75518
rect 25116 75572 25172 79200
rect 25788 76580 25844 79200
rect 26124 76580 26180 76590
rect 25788 76578 26180 76580
rect 25788 76526 26126 76578
rect 26178 76526 26180 76578
rect 25788 76524 26180 76526
rect 26124 76514 26180 76524
rect 26796 76580 26852 76590
rect 26796 75794 26852 76524
rect 26796 75742 26798 75794
rect 26850 75742 26852 75794
rect 26796 75730 26852 75742
rect 25340 75572 25396 75582
rect 25116 75570 25396 75572
rect 25116 75518 25342 75570
rect 25394 75518 25396 75570
rect 25116 75516 25396 75518
rect 27132 75572 27188 79200
rect 27244 76580 27300 76590
rect 27244 76466 27300 76524
rect 27244 76414 27246 76466
rect 27298 76414 27300 76466
rect 27244 76402 27300 76414
rect 27804 76356 27860 79200
rect 29148 77252 29204 79200
rect 28700 77196 29204 77252
rect 27804 76290 27860 76300
rect 28252 76466 28308 76478
rect 28252 76414 28254 76466
rect 28306 76414 28308 76466
rect 27356 75572 27412 75582
rect 27132 75570 27412 75572
rect 27132 75518 27358 75570
rect 27410 75518 27412 75570
rect 27132 75516 27412 75518
rect 21756 75478 21812 75516
rect 23324 75506 23380 75516
rect 25340 75506 25396 75516
rect 27356 75506 27412 75516
rect 28252 75570 28308 76414
rect 28252 75518 28254 75570
rect 28306 75518 28308 75570
rect 28252 75506 28308 75518
rect 28588 75570 28644 75582
rect 28588 75518 28590 75570
rect 28642 75518 28644 75570
rect 21644 74946 21700 74956
rect 28588 74340 28644 75518
rect 28700 75122 28756 77196
rect 29260 76468 29316 76478
rect 28812 76356 28868 76366
rect 28812 76262 28868 76300
rect 29260 75572 29316 76412
rect 29820 76356 29876 79200
rect 30044 76468 30100 76478
rect 29820 76290 29876 76300
rect 29932 76466 30100 76468
rect 29932 76414 30046 76466
rect 30098 76414 30100 76466
rect 29932 76412 30100 76414
rect 29484 76020 29540 76030
rect 29484 75906 29540 75964
rect 29484 75854 29486 75906
rect 29538 75854 29540 75906
rect 29484 75842 29540 75854
rect 29372 75796 29428 75806
rect 29372 75702 29428 75740
rect 28700 75070 28702 75122
rect 28754 75070 28756 75122
rect 28700 75058 28756 75070
rect 29148 75570 29316 75572
rect 29148 75518 29262 75570
rect 29314 75518 29316 75570
rect 29148 75516 29316 75518
rect 28588 74274 28644 74284
rect 28924 74788 28980 74798
rect 28924 74226 28980 74732
rect 28924 74174 28926 74226
rect 28978 74174 28980 74226
rect 28924 74162 28980 74174
rect 29148 73892 29204 75516
rect 29260 75506 29316 75516
rect 29932 75236 29988 76412
rect 30044 76402 30100 76412
rect 30716 76356 30772 76366
rect 30716 76262 30772 76300
rect 31164 76132 31220 79200
rect 31836 76356 31892 79200
rect 33180 77812 33236 79200
rect 33180 77756 33460 77812
rect 33180 77588 33236 77598
rect 33068 76580 33124 76590
rect 31836 76290 31892 76300
rect 32172 76466 32228 76478
rect 32172 76414 32174 76466
rect 32226 76414 32228 76466
rect 31164 76076 31556 76132
rect 30828 75796 30884 75806
rect 30044 75684 30100 75694
rect 30044 75590 30100 75628
rect 30380 75682 30436 75694
rect 30380 75630 30382 75682
rect 30434 75630 30436 75682
rect 29372 75180 29988 75236
rect 30268 75572 30324 75582
rect 29372 75122 29428 75180
rect 29372 75070 29374 75122
rect 29426 75070 29428 75122
rect 29372 75058 29428 75070
rect 30268 75122 30324 75516
rect 30268 75070 30270 75122
rect 30322 75070 30324 75122
rect 30268 75058 30324 75070
rect 29932 75012 29988 75022
rect 29932 74918 29988 74956
rect 29372 74900 29428 74910
rect 29260 74788 29316 74798
rect 29260 74694 29316 74732
rect 29260 74228 29316 74238
rect 29372 74228 29428 74844
rect 29260 74226 29428 74228
rect 29260 74174 29262 74226
rect 29314 74174 29428 74226
rect 29260 74172 29428 74174
rect 29820 74228 29876 74238
rect 29260 74162 29316 74172
rect 29820 74134 29876 74172
rect 29148 73826 29204 73836
rect 30268 73892 30324 73902
rect 30268 73798 30324 73836
rect 19836 73724 20100 73734
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 19836 73658 20100 73668
rect 30380 73218 30436 75630
rect 30492 75684 30548 75694
rect 30492 74114 30548 75628
rect 30604 75682 30660 75694
rect 30604 75630 30606 75682
rect 30658 75630 30660 75682
rect 30604 75572 30660 75630
rect 30604 75506 30660 75516
rect 30828 75010 30884 75740
rect 31164 75682 31220 75694
rect 31164 75630 31166 75682
rect 31218 75630 31220 75682
rect 31164 75572 31220 75630
rect 31164 75506 31220 75516
rect 31388 75682 31444 75694
rect 31388 75630 31390 75682
rect 31442 75630 31444 75682
rect 31276 75460 31332 75470
rect 31276 75122 31332 75404
rect 31388 75236 31444 75630
rect 31388 75170 31444 75180
rect 31276 75070 31278 75122
rect 31330 75070 31332 75122
rect 31276 75058 31332 75070
rect 30828 74958 30830 75010
rect 30882 74958 30884 75010
rect 30828 74946 30884 74958
rect 31164 75012 31220 75022
rect 31052 74898 31108 74910
rect 31052 74846 31054 74898
rect 31106 74846 31108 74898
rect 31052 74228 31108 74846
rect 31052 74162 31108 74172
rect 30492 74062 30494 74114
rect 30546 74062 30548 74114
rect 30492 74050 30548 74062
rect 31164 74114 31220 74956
rect 31388 74900 31444 74910
rect 31164 74062 31166 74114
rect 31218 74062 31220 74114
rect 31164 73892 31220 74062
rect 30940 73836 31220 73892
rect 31276 74898 31444 74900
rect 31276 74846 31390 74898
rect 31442 74846 31444 74898
rect 31276 74844 31444 74846
rect 30940 73554 30996 73836
rect 30940 73502 30942 73554
rect 30994 73502 30996 73554
rect 30940 73490 30996 73502
rect 30380 73166 30382 73218
rect 30434 73166 30436 73218
rect 30380 72660 30436 73166
rect 30380 72594 30436 72604
rect 31276 72660 31332 74844
rect 31388 74834 31444 74844
rect 31500 74676 31556 76076
rect 32172 76020 32228 76414
rect 32732 76356 32788 76366
rect 32732 76262 32788 76300
rect 31724 75684 31780 75694
rect 31724 75682 32004 75684
rect 31724 75630 31726 75682
rect 31778 75630 32004 75682
rect 31724 75628 32004 75630
rect 31724 75618 31780 75628
rect 31388 74620 31556 74676
rect 31836 75236 31892 75246
rect 31388 73554 31444 74620
rect 31836 74228 31892 75180
rect 31836 74004 31892 74172
rect 31948 74116 32004 75628
rect 32060 75572 32116 75582
rect 32060 74900 32116 75516
rect 32172 75236 32228 75964
rect 32284 75572 32340 75582
rect 32620 75572 32676 75582
rect 32284 75570 32564 75572
rect 32284 75518 32286 75570
rect 32338 75518 32564 75570
rect 32284 75516 32564 75518
rect 32284 75506 32340 75516
rect 32508 75236 32564 75516
rect 32620 75478 32676 75516
rect 32172 75180 32452 75236
rect 32060 74768 32116 74844
rect 32284 74788 32340 74798
rect 32060 74116 32116 74126
rect 31948 74114 32116 74116
rect 31948 74062 32062 74114
rect 32114 74062 32116 74114
rect 31948 74060 32116 74062
rect 32060 74050 32116 74060
rect 31836 73948 32004 74004
rect 31500 73892 31556 73902
rect 31500 73798 31556 73836
rect 31388 73502 31390 73554
rect 31442 73502 31444 73554
rect 31388 73490 31444 73502
rect 31948 72996 32004 73948
rect 32172 73556 32228 73566
rect 32284 73556 32340 74732
rect 32396 74002 32452 75180
rect 32508 75170 32564 75180
rect 33068 74788 33124 76524
rect 33180 75570 33236 77532
rect 33180 75518 33182 75570
rect 33234 75518 33236 75570
rect 33180 75460 33236 75518
rect 33180 75394 33236 75404
rect 33292 75458 33348 75470
rect 33292 75406 33294 75458
rect 33346 75406 33348 75458
rect 33180 75236 33236 75246
rect 33180 75122 33236 75180
rect 33180 75070 33182 75122
rect 33234 75070 33236 75122
rect 33180 75058 33236 75070
rect 33292 75124 33348 75406
rect 33292 75058 33348 75068
rect 33068 74732 33236 74788
rect 32620 74676 32676 74686
rect 32620 74674 33124 74676
rect 32620 74622 32622 74674
rect 32674 74622 33124 74674
rect 32620 74620 33124 74622
rect 32620 74610 32676 74620
rect 32396 73950 32398 74002
rect 32450 73950 32452 74002
rect 32396 73938 32452 73950
rect 32732 74116 32788 74126
rect 32172 73554 32676 73556
rect 32172 73502 32174 73554
rect 32226 73502 32676 73554
rect 32172 73500 32676 73502
rect 32172 73490 32228 73500
rect 32620 73332 32676 73500
rect 32732 73554 32788 74060
rect 33068 74114 33124 74620
rect 33068 74062 33070 74114
rect 33122 74062 33124 74114
rect 33068 74050 33124 74062
rect 33180 73892 33236 74732
rect 33404 74116 33460 77756
rect 33852 77250 33908 79200
rect 33852 77198 33854 77250
rect 33906 77198 33908 77250
rect 33852 77186 33908 77198
rect 34748 77250 34804 77262
rect 34748 77198 34750 77250
rect 34802 77198 34804 77250
rect 34076 76466 34132 76478
rect 34076 76414 34078 76466
rect 34130 76414 34132 76466
rect 33516 75570 33572 75582
rect 33740 75572 33796 75582
rect 33516 75518 33518 75570
rect 33570 75518 33572 75570
rect 33516 74676 33572 75518
rect 33516 74582 33572 74620
rect 33628 75570 33796 75572
rect 33628 75518 33742 75570
rect 33794 75518 33796 75570
rect 33628 75516 33796 75518
rect 33628 74340 33684 75516
rect 33740 75506 33796 75516
rect 33852 75572 33908 75582
rect 33740 74900 33796 74910
rect 33740 74806 33796 74844
rect 33404 74050 33460 74060
rect 33516 74284 33684 74340
rect 33404 73892 33460 73902
rect 33180 73890 33460 73892
rect 33180 73838 33406 73890
rect 33458 73838 33460 73890
rect 33180 73836 33460 73838
rect 32732 73502 32734 73554
rect 32786 73502 32788 73554
rect 32732 73490 32788 73502
rect 32620 73276 32900 73332
rect 31948 72940 32452 72996
rect 31276 72594 31332 72604
rect 31836 72660 31892 72670
rect 15820 72258 15876 72268
rect 19836 72156 20100 72166
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 19836 72090 20100 72100
rect 13804 71474 13860 71484
rect 4476 71372 4740 71382
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4476 71306 4740 71316
rect 19836 70588 20100 70598
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 19836 70522 20100 70532
rect 31836 70420 31892 72604
rect 31948 72660 32004 72670
rect 31948 72566 32004 72604
rect 32396 72658 32452 72940
rect 32396 72606 32398 72658
rect 32450 72606 32452 72658
rect 32396 72594 32452 72606
rect 32844 72658 32900 73276
rect 32844 72606 32846 72658
rect 32898 72606 32900 72658
rect 32844 72594 32900 72606
rect 33292 72658 33348 73836
rect 33404 73554 33460 73836
rect 33404 73502 33406 73554
rect 33458 73502 33460 73554
rect 33404 73490 33460 73502
rect 33516 73554 33572 74284
rect 33852 73892 33908 75516
rect 34076 75572 34132 76414
rect 34636 76468 34692 76478
rect 34076 75506 34132 75516
rect 34412 75572 34468 75582
rect 34412 75478 34468 75516
rect 34300 75460 34356 75470
rect 33964 74340 34020 74350
rect 33964 74246 34020 74284
rect 34300 74338 34356 75404
rect 34636 75122 34692 76412
rect 34748 76354 34804 77198
rect 35196 76468 35252 79200
rect 35868 77812 35924 79200
rect 35868 77756 36820 77812
rect 34748 76302 34750 76354
rect 34802 76302 34804 76354
rect 34748 76290 34804 76302
rect 34860 76412 35252 76468
rect 35756 77252 35812 77262
rect 34636 75070 34638 75122
rect 34690 75070 34692 75122
rect 34636 75058 34692 75070
rect 34300 74286 34302 74338
rect 34354 74286 34356 74338
rect 33516 73502 33518 73554
rect 33570 73502 33572 73554
rect 33516 73490 33572 73502
rect 33628 73836 33908 73892
rect 33628 73442 33684 73836
rect 34188 73780 34244 73790
rect 34188 73444 34244 73724
rect 33628 73390 33630 73442
rect 33682 73390 33684 73442
rect 33628 73378 33684 73390
rect 33852 73442 34244 73444
rect 33852 73390 34190 73442
rect 34242 73390 34244 73442
rect 33852 73388 34244 73390
rect 33292 72606 33294 72658
rect 33346 72606 33348 72658
rect 33292 72594 33348 72606
rect 33740 72770 33796 72782
rect 33740 72718 33742 72770
rect 33794 72718 33796 72770
rect 33740 72658 33796 72718
rect 33740 72606 33742 72658
rect 33794 72606 33796 72658
rect 33740 72594 33796 72606
rect 33852 71986 33908 73388
rect 34188 73378 34244 73388
rect 34300 72770 34356 74286
rect 34412 74898 34468 74910
rect 34412 74846 34414 74898
rect 34466 74846 34468 74898
rect 34412 74340 34468 74846
rect 34412 74274 34468 74284
rect 34524 74228 34580 74238
rect 34524 73554 34580 74172
rect 34524 73502 34526 73554
rect 34578 73502 34580 73554
rect 34524 73490 34580 73502
rect 34300 72718 34302 72770
rect 34354 72718 34356 72770
rect 34188 72660 34244 72670
rect 34188 72566 34244 72604
rect 33852 71934 33854 71986
rect 33906 71934 33908 71986
rect 33852 71922 33908 71934
rect 34300 71092 34356 72718
rect 34748 72436 34804 72446
rect 34860 72436 34916 76412
rect 35084 76244 35140 76254
rect 35084 75794 35140 76188
rect 35196 76076 35460 76086
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35196 76010 35460 76020
rect 35084 75742 35086 75794
rect 35138 75742 35140 75794
rect 35084 75730 35140 75742
rect 34972 75570 35028 75582
rect 34972 75518 34974 75570
rect 35026 75518 35028 75570
rect 34972 75460 35028 75518
rect 34972 75394 35028 75404
rect 35308 75570 35364 75582
rect 35308 75518 35310 75570
rect 35362 75518 35364 75570
rect 35196 74900 35252 74910
rect 35308 74900 35364 75518
rect 35532 75570 35588 75582
rect 35532 75518 35534 75570
rect 35586 75518 35588 75570
rect 35532 75124 35588 75518
rect 35756 75460 35812 77196
rect 36092 76468 36148 76478
rect 36092 76374 36148 76412
rect 36764 76354 36820 77756
rect 36764 76302 36766 76354
rect 36818 76302 36820 76354
rect 36764 76290 36820 76302
rect 35644 75124 35700 75134
rect 35532 75122 35700 75124
rect 35532 75070 35646 75122
rect 35698 75070 35700 75122
rect 35532 75068 35700 75070
rect 35644 75058 35700 75068
rect 35756 75122 35812 75404
rect 35756 75070 35758 75122
rect 35810 75070 35812 75122
rect 35756 75058 35812 75070
rect 35980 76244 36036 76254
rect 35532 74900 35588 74910
rect 35308 74898 35588 74900
rect 35308 74846 35534 74898
rect 35586 74846 35588 74898
rect 35308 74844 35588 74846
rect 35196 74806 35252 74844
rect 35532 74788 35588 74844
rect 35196 74508 35460 74518
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35196 74442 35460 74452
rect 35084 74340 35140 74350
rect 35084 74246 35140 74284
rect 35420 74340 35476 74350
rect 35532 74340 35588 74732
rect 35420 74338 35588 74340
rect 35420 74286 35422 74338
rect 35474 74286 35588 74338
rect 35420 74284 35588 74286
rect 35644 74900 35700 74910
rect 35420 74274 35476 74284
rect 35644 74228 35700 74844
rect 35308 74116 35364 74126
rect 35644 74096 35700 74172
rect 35756 74452 35812 74462
rect 35308 73442 35364 74060
rect 35756 74004 35812 74396
rect 35420 73948 35812 74004
rect 35420 73554 35476 73948
rect 35420 73502 35422 73554
rect 35474 73502 35476 73554
rect 35420 73490 35476 73502
rect 35308 73390 35310 73442
rect 35362 73390 35364 73442
rect 35308 73378 35364 73390
rect 35980 73442 36036 76188
rect 36652 76132 36708 76142
rect 36316 75908 36372 75918
rect 36316 75794 36372 75852
rect 36316 75742 36318 75794
rect 36370 75742 36372 75794
rect 36316 75730 36372 75742
rect 36652 75572 36708 76076
rect 36540 75570 36708 75572
rect 36540 75518 36654 75570
rect 36706 75518 36708 75570
rect 36540 75516 36708 75518
rect 36316 75460 36372 75470
rect 36204 75458 36372 75460
rect 36204 75406 36318 75458
rect 36370 75406 36372 75458
rect 36204 75404 36372 75406
rect 35980 73390 35982 73442
rect 36034 73390 36036 73442
rect 35532 73108 35588 73118
rect 35196 72940 35460 72950
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35196 72874 35460 72884
rect 35420 72660 35476 72670
rect 35532 72660 35588 73052
rect 35476 72604 35588 72660
rect 35420 72528 35476 72604
rect 34748 72434 34916 72436
rect 34748 72382 34750 72434
rect 34802 72382 34916 72434
rect 34748 72380 34916 72382
rect 34748 72370 34804 72380
rect 35308 72324 35364 72334
rect 35308 72230 35364 72268
rect 35980 71986 36036 73390
rect 35980 71934 35982 71986
rect 36034 71934 36036 71986
rect 35980 71922 36036 71934
rect 36092 73442 36148 73454
rect 36092 73390 36094 73442
rect 36146 73390 36148 73442
rect 34972 71652 35028 71662
rect 35420 71652 35476 71662
rect 34972 71650 35588 71652
rect 34972 71598 34974 71650
rect 35026 71598 35422 71650
rect 35474 71598 35588 71650
rect 34972 71596 35588 71598
rect 34972 71586 35028 71596
rect 35420 71586 35476 71596
rect 34860 71540 34916 71550
rect 34860 71446 34916 71484
rect 35196 71372 35460 71382
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35196 71306 35460 71316
rect 34300 71026 34356 71036
rect 35196 71092 35252 71102
rect 35196 70998 35252 71036
rect 35532 70532 35588 71596
rect 35644 71092 35700 71102
rect 35644 70998 35700 71036
rect 36092 70980 36148 73390
rect 36092 70914 36148 70924
rect 36204 71316 36260 75404
rect 36316 75394 36372 75404
rect 36428 75458 36484 75470
rect 36428 75406 36430 75458
rect 36482 75406 36484 75458
rect 36428 75122 36484 75406
rect 36428 75070 36430 75122
rect 36482 75070 36484 75122
rect 36428 75058 36484 75070
rect 36540 75012 36596 75516
rect 36652 75506 36708 75516
rect 36876 75570 36932 75582
rect 36876 75518 36878 75570
rect 36930 75518 36932 75570
rect 36316 74676 36372 74686
rect 36316 74338 36372 74620
rect 36316 74286 36318 74338
rect 36370 74286 36372 74338
rect 36316 74274 36372 74286
rect 36316 74004 36372 74014
rect 36316 73554 36372 73948
rect 36316 73502 36318 73554
rect 36370 73502 36372 73554
rect 36316 73490 36372 73502
rect 36428 72436 36484 72446
rect 36428 72342 36484 72380
rect 36428 71988 36484 71998
rect 36428 71894 36484 71932
rect 36092 70756 36148 70766
rect 36204 70756 36260 71260
rect 36428 70980 36484 70990
rect 36428 70886 36484 70924
rect 36092 70754 36260 70756
rect 36092 70702 36094 70754
rect 36146 70702 36260 70754
rect 36092 70700 36260 70702
rect 36092 70690 36148 70700
rect 35532 70466 35588 70476
rect 31836 70354 31892 70364
rect 36540 70196 36596 74956
rect 36876 74788 36932 75518
rect 37212 74788 37268 79200
rect 37884 76804 37940 79200
rect 37884 76738 37940 76748
rect 38332 76692 38388 76702
rect 37884 76578 37940 76590
rect 37884 76526 37886 76578
rect 37938 76526 37940 76578
rect 37548 75460 37604 75470
rect 37548 75366 37604 75404
rect 37548 75236 37604 75246
rect 37324 75012 37380 75022
rect 37324 74918 37380 74956
rect 37548 74900 37604 75180
rect 37884 75236 37940 76526
rect 38108 76468 38164 76478
rect 37884 75170 37940 75180
rect 37996 76466 38164 76468
rect 37996 76414 38110 76466
rect 38162 76414 38164 76466
rect 37996 76412 38164 76414
rect 37996 76020 38052 76412
rect 38108 76402 38164 76412
rect 37436 74898 37604 74900
rect 37436 74846 37550 74898
rect 37602 74846 37604 74898
rect 37436 74844 37604 74846
rect 37212 74732 37380 74788
rect 36764 74674 36820 74686
rect 36764 74622 36766 74674
rect 36818 74622 36820 74674
rect 36652 74114 36708 74126
rect 36652 74062 36654 74114
rect 36706 74062 36708 74114
rect 36652 73554 36708 74062
rect 36652 73502 36654 73554
rect 36706 73502 36708 73554
rect 36652 73490 36708 73502
rect 36764 70420 36820 74622
rect 36876 74228 36932 74732
rect 36876 74162 36932 74172
rect 37212 74002 37268 74014
rect 37212 73950 37214 74002
rect 37266 73950 37268 74002
rect 36876 73556 36932 73566
rect 36876 73462 36932 73500
rect 36988 73330 37044 73342
rect 36988 73278 36990 73330
rect 37042 73278 37044 73330
rect 36988 72996 37044 73278
rect 36988 72930 37044 72940
rect 37212 72772 37268 73950
rect 36988 72716 37268 72772
rect 36988 72658 37044 72716
rect 36988 72606 36990 72658
rect 37042 72606 37044 72658
rect 36988 72594 37044 72606
rect 37324 72324 37380 74732
rect 37436 74114 37492 74844
rect 37548 74834 37604 74844
rect 37436 74062 37438 74114
rect 37490 74062 37492 74114
rect 37436 74050 37492 74062
rect 37548 73668 37604 73678
rect 37548 73442 37604 73612
rect 37548 73390 37550 73442
rect 37602 73390 37604 73442
rect 37548 73378 37604 73390
rect 37772 73668 37828 73678
rect 37660 73332 37716 73342
rect 37548 72996 37604 73006
rect 36988 72268 37380 72324
rect 37436 72660 37492 72670
rect 37436 72546 37492 72604
rect 37436 72494 37438 72546
rect 37490 72494 37492 72546
rect 36988 71986 37044 72268
rect 37436 72212 37492 72494
rect 36988 71934 36990 71986
rect 37042 71934 37044 71986
rect 36988 71922 37044 71934
rect 37324 72156 37492 72212
rect 37324 71090 37380 72156
rect 37436 71988 37492 71998
rect 37548 71988 37604 72940
rect 37436 71986 37604 71988
rect 37436 71934 37438 71986
rect 37490 71934 37604 71986
rect 37436 71932 37604 71934
rect 37660 71986 37716 73276
rect 37660 71934 37662 71986
rect 37714 71934 37716 71986
rect 37436 71922 37492 71932
rect 37660 71922 37716 71934
rect 37772 71988 37828 73612
rect 37884 73444 37940 73454
rect 37884 73350 37940 73388
rect 37884 72548 37940 72558
rect 37884 72454 37940 72492
rect 37772 71874 37828 71932
rect 37772 71822 37774 71874
rect 37826 71822 37828 71874
rect 37324 71038 37326 71090
rect 37378 71038 37380 71090
rect 37324 71026 37380 71038
rect 37660 71092 37716 71102
rect 37772 71092 37828 71822
rect 37660 71090 37828 71092
rect 37660 71038 37662 71090
rect 37714 71038 37828 71090
rect 37660 71036 37828 71038
rect 37660 71026 37716 71036
rect 37772 70868 37828 71036
rect 37772 70802 37828 70812
rect 36764 70354 36820 70364
rect 36540 70130 36596 70140
rect 37212 70196 37268 70206
rect 37212 70102 37268 70140
rect 37548 70196 37604 70206
rect 37548 70102 37604 70140
rect 37996 69970 38052 75964
rect 38108 75682 38164 75694
rect 38108 75630 38110 75682
rect 38162 75630 38164 75682
rect 38108 74452 38164 75630
rect 38220 74900 38276 74910
rect 38220 74806 38276 74844
rect 38108 74386 38164 74396
rect 38220 74340 38276 74350
rect 38332 74340 38388 76636
rect 38556 76580 38612 79200
rect 38556 76514 38612 76524
rect 38780 76804 38836 76814
rect 38780 75794 38836 76748
rect 39116 76580 39172 76590
rect 38780 75742 38782 75794
rect 38834 75742 38836 75794
rect 38780 75730 38836 75742
rect 38892 75908 38948 75918
rect 38668 75684 38724 75694
rect 38220 74338 38388 74340
rect 38220 74286 38222 74338
rect 38274 74286 38388 74338
rect 38220 74284 38388 74286
rect 38556 75012 38612 75022
rect 38220 74274 38276 74284
rect 38108 74116 38164 74126
rect 38108 70980 38164 74060
rect 38556 74004 38612 74956
rect 38668 75010 38724 75628
rect 38780 75460 38836 75470
rect 38780 75236 38836 75404
rect 38780 75122 38836 75180
rect 38780 75070 38782 75122
rect 38834 75070 38836 75122
rect 38780 75058 38836 75070
rect 38668 74958 38670 75010
rect 38722 74958 38724 75010
rect 38668 74946 38724 74958
rect 38668 74788 38724 74798
rect 38668 74694 38724 74732
rect 38780 74116 38836 74126
rect 38892 74116 38948 75852
rect 39004 75012 39060 75022
rect 39004 74918 39060 74956
rect 38780 74114 38948 74116
rect 38780 74062 38782 74114
rect 38834 74062 38948 74114
rect 38780 74060 38948 74062
rect 38556 73948 38724 74004
rect 38444 73892 38500 73902
rect 38444 73332 38500 73836
rect 38668 73332 38724 73948
rect 38780 73668 38836 74060
rect 38780 73602 38836 73612
rect 38892 73890 38948 73902
rect 38892 73838 38894 73890
rect 38946 73838 38948 73890
rect 38892 73556 38948 73838
rect 39004 73892 39060 73902
rect 39004 73798 39060 73836
rect 38892 73490 38948 73500
rect 38892 73332 38948 73342
rect 38500 73276 38612 73332
rect 38668 73276 38836 73332
rect 38444 73200 38500 73276
rect 38444 72548 38500 72558
rect 38556 72548 38612 73276
rect 38668 73106 38724 73118
rect 38668 73054 38670 73106
rect 38722 73054 38724 73106
rect 38668 72884 38724 73054
rect 38668 72818 38724 72828
rect 38556 72492 38724 72548
rect 38444 71986 38500 72492
rect 38556 72324 38612 72334
rect 38556 72230 38612 72268
rect 38444 71934 38446 71986
rect 38498 71934 38500 71986
rect 38444 71922 38500 71934
rect 38220 71092 38276 71102
rect 38220 70998 38276 71036
rect 38108 70418 38164 70924
rect 38668 70866 38724 72492
rect 38780 71988 38836 73276
rect 38780 71922 38836 71932
rect 38668 70814 38670 70866
rect 38722 70814 38724 70866
rect 38668 70802 38724 70814
rect 38780 71764 38836 71774
rect 38780 70532 38836 71708
rect 38892 70644 38948 73276
rect 39004 73106 39060 73118
rect 39004 73054 39006 73106
rect 39058 73054 39060 73106
rect 39004 72546 39060 73054
rect 39004 72494 39006 72546
rect 39058 72494 39060 72546
rect 39004 72482 39060 72494
rect 39004 72324 39060 72334
rect 39004 71764 39060 72268
rect 39004 71698 39060 71708
rect 39004 71540 39060 71550
rect 39004 71092 39060 71484
rect 39004 70978 39060 71036
rect 39004 70926 39006 70978
rect 39058 70926 39060 70978
rect 39004 70914 39060 70926
rect 39004 70644 39060 70654
rect 38892 70588 39004 70644
rect 38108 70366 38110 70418
rect 38162 70366 38164 70418
rect 38108 70354 38164 70366
rect 38556 70476 38836 70532
rect 38556 70418 38612 70476
rect 38556 70366 38558 70418
rect 38610 70366 38612 70418
rect 38556 70354 38612 70366
rect 39004 70418 39060 70588
rect 39004 70366 39006 70418
rect 39058 70366 39060 70418
rect 39004 70354 39060 70366
rect 37996 69918 37998 69970
rect 38050 69918 38052 69970
rect 37996 69906 38052 69918
rect 38556 69970 38612 69982
rect 38556 69918 38558 69970
rect 38610 69918 38612 69970
rect 4476 69804 4740 69814
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4476 69738 4740 69748
rect 35196 69804 35460 69814
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35196 69738 35460 69748
rect 38556 69522 38612 69918
rect 38556 69470 38558 69522
rect 38610 69470 38612 69522
rect 38556 69458 38612 69470
rect 39004 69524 39060 69534
rect 39116 69524 39172 76524
rect 39228 72436 39284 79200
rect 39228 72370 39284 72380
rect 39340 76356 39396 76366
rect 39340 74114 39396 76300
rect 39900 75796 39956 79200
rect 40572 77026 40628 79200
rect 40572 76974 40574 77026
rect 40626 76974 40628 77026
rect 40572 76962 40628 76974
rect 40908 76692 40964 76702
rect 41244 76692 41300 79200
rect 40908 76690 41300 76692
rect 40908 76638 40910 76690
rect 40962 76638 41300 76690
rect 40908 76636 41300 76638
rect 41804 77026 41860 77038
rect 41804 76974 41806 77026
rect 41858 76974 41860 77026
rect 40908 76626 40964 76636
rect 40012 76354 40068 76366
rect 40012 76302 40014 76354
rect 40066 76302 40068 76354
rect 40012 76244 40068 76302
rect 41692 76356 41748 76366
rect 41692 76262 41748 76300
rect 40012 76178 40068 76188
rect 39900 75730 39956 75740
rect 40236 75908 40292 75918
rect 40236 75684 40292 75852
rect 40460 75796 40516 75806
rect 40460 75702 40516 75740
rect 40236 75628 40404 75684
rect 40012 75572 40068 75582
rect 39676 75570 40068 75572
rect 39676 75518 40014 75570
rect 40066 75518 40068 75570
rect 39676 75516 40068 75518
rect 39676 75460 39732 75516
rect 40012 75506 40068 75516
rect 39340 74062 39342 74114
rect 39394 74062 39396 74114
rect 39228 71988 39284 71998
rect 39228 70980 39284 71932
rect 39228 70196 39284 70924
rect 39228 70130 39284 70140
rect 39340 69860 39396 74062
rect 39452 75404 39732 75460
rect 40124 75458 40180 75470
rect 40124 75406 40126 75458
rect 40178 75406 40180 75458
rect 39452 74898 39508 75404
rect 40124 75348 40180 75406
rect 40124 75282 40180 75292
rect 40236 75458 40292 75470
rect 40236 75406 40238 75458
rect 40290 75406 40292 75458
rect 40012 75124 40068 75134
rect 40012 75030 40068 75068
rect 40124 75124 40180 75134
rect 40236 75124 40292 75406
rect 40124 75122 40292 75124
rect 40124 75070 40126 75122
rect 40178 75070 40292 75122
rect 40124 75068 40292 75070
rect 40124 75058 40180 75068
rect 40236 75012 40292 75068
rect 40236 74946 40292 74956
rect 39452 74846 39454 74898
rect 39506 74846 39508 74898
rect 39452 74004 39508 74846
rect 39900 74898 39956 74910
rect 39900 74846 39902 74898
rect 39954 74846 39956 74898
rect 39900 74788 39956 74846
rect 40348 74788 40404 75628
rect 40684 75682 40740 75694
rect 40684 75630 40686 75682
rect 40738 75630 40740 75682
rect 39900 74732 40404 74788
rect 40460 75572 40516 75582
rect 40012 74228 40068 74238
rect 39452 73938 39508 73948
rect 39900 74004 39956 74042
rect 39900 73938 39956 73948
rect 39676 73892 39732 73902
rect 39676 73554 39732 73836
rect 39676 73502 39678 73554
rect 39730 73502 39732 73554
rect 39676 73490 39732 73502
rect 40012 73332 40068 74172
rect 40348 74228 40404 74238
rect 40348 74114 40404 74172
rect 40348 74062 40350 74114
rect 40402 74062 40404 74114
rect 40348 74050 40404 74062
rect 40460 74226 40516 75516
rect 40684 75124 40740 75630
rect 41132 75684 41188 75694
rect 41132 75590 41188 75628
rect 41692 75572 41748 75582
rect 41692 75478 41748 75516
rect 41244 75460 41300 75470
rect 41468 75460 41524 75470
rect 41244 75366 41300 75404
rect 41356 75458 41524 75460
rect 41356 75406 41470 75458
rect 41522 75406 41524 75458
rect 41356 75404 41524 75406
rect 41132 75348 41188 75358
rect 40684 75058 40740 75068
rect 41020 75124 41076 75134
rect 41020 75030 41076 75068
rect 40796 75012 40852 75022
rect 40796 74898 40852 74956
rect 40796 74846 40798 74898
rect 40850 74846 40852 74898
rect 40796 74834 40852 74846
rect 40908 74900 40964 74910
rect 40460 74174 40462 74226
rect 40514 74174 40516 74226
rect 40012 73266 40068 73276
rect 39788 73218 39844 73230
rect 39788 73166 39790 73218
rect 39842 73166 39844 73218
rect 39676 72546 39732 72558
rect 39676 72494 39678 72546
rect 39730 72494 39732 72546
rect 39676 71876 39732 72494
rect 39788 72548 39844 73166
rect 39900 73108 39956 73118
rect 39900 73106 40068 73108
rect 39900 73054 39902 73106
rect 39954 73054 40068 73106
rect 39900 73052 40068 73054
rect 39900 73042 39956 73052
rect 40012 72884 40068 73052
rect 39900 72548 39956 72558
rect 39788 72546 39956 72548
rect 39788 72494 39902 72546
rect 39954 72494 39956 72546
rect 39788 72492 39956 72494
rect 39900 72482 39956 72492
rect 40012 72324 40068 72828
rect 40348 72548 40404 72558
rect 40348 72454 40404 72492
rect 40012 72258 40068 72268
rect 40236 72434 40292 72446
rect 40236 72382 40238 72434
rect 40290 72382 40292 72434
rect 40124 71876 40180 71886
rect 39676 71820 39844 71876
rect 39788 71762 39844 71820
rect 39788 71710 39790 71762
rect 39842 71710 39844 71762
rect 39788 71204 39844 71710
rect 40124 71540 40180 71820
rect 40124 71474 40180 71484
rect 39452 71148 39844 71204
rect 39900 71204 39956 71214
rect 39452 70418 39508 71148
rect 39900 71110 39956 71148
rect 40236 71092 40292 72382
rect 40236 71026 40292 71036
rect 40348 71204 40404 71214
rect 39452 70366 39454 70418
rect 39506 70366 39508 70418
rect 39452 70354 39508 70366
rect 39676 70868 39732 70878
rect 39564 70082 39620 70094
rect 39564 70030 39566 70082
rect 39618 70030 39620 70082
rect 39564 69860 39620 70030
rect 39340 69804 39620 69860
rect 39004 69522 39172 69524
rect 39004 69470 39006 69522
rect 39058 69470 39172 69522
rect 39004 69468 39172 69470
rect 39676 69522 39732 70812
rect 39788 70866 39844 70878
rect 39788 70814 39790 70866
rect 39842 70814 39844 70866
rect 39788 70644 39844 70814
rect 39900 70756 39956 70766
rect 39900 70662 39956 70700
rect 39788 70578 39844 70588
rect 40124 70420 40180 70430
rect 40124 70326 40180 70364
rect 40348 70418 40404 71148
rect 40348 70366 40350 70418
rect 40402 70366 40404 70418
rect 40348 70354 40404 70366
rect 40460 70306 40516 74174
rect 40572 74002 40628 74014
rect 40572 73950 40574 74002
rect 40626 73950 40628 74002
rect 40572 73892 40628 73950
rect 40796 74004 40852 74042
rect 40796 73938 40852 73948
rect 40572 73826 40628 73836
rect 40908 73554 40964 74844
rect 40908 73502 40910 73554
rect 40962 73502 40964 73554
rect 40908 73490 40964 73502
rect 41020 74004 41076 74014
rect 41020 73556 41076 73948
rect 41020 73490 41076 73500
rect 40572 73442 40628 73454
rect 40572 73390 40574 73442
rect 40626 73390 40628 73442
rect 40572 73220 40628 73390
rect 40796 73332 40852 73342
rect 40796 73238 40852 73276
rect 41020 73330 41076 73342
rect 41020 73278 41022 73330
rect 41074 73278 41076 73330
rect 40572 73154 40628 73164
rect 41020 73108 41076 73278
rect 41020 73042 41076 73052
rect 41020 72772 41076 72782
rect 40572 72660 40628 72670
rect 40572 72546 40628 72604
rect 40572 72494 40574 72546
rect 40626 72494 40628 72546
rect 40572 72482 40628 72494
rect 41020 71986 41076 72716
rect 41132 72660 41188 75292
rect 41356 73948 41412 75404
rect 41468 75394 41524 75404
rect 41692 74788 41748 74798
rect 41132 72594 41188 72604
rect 41244 73892 41412 73948
rect 41468 74786 41748 74788
rect 41468 74734 41694 74786
rect 41746 74734 41748 74786
rect 41468 74732 41748 74734
rect 41468 73892 41524 74732
rect 41692 74722 41748 74732
rect 41692 74114 41748 74126
rect 41692 74062 41694 74114
rect 41746 74062 41748 74114
rect 41692 73948 41748 74062
rect 41020 71934 41022 71986
rect 41074 71934 41076 71986
rect 41020 71876 41076 71934
rect 41020 71810 41076 71820
rect 41132 71652 41188 71662
rect 40908 71092 40964 71102
rect 40908 70998 40964 71036
rect 41132 70978 41188 71596
rect 41244 71204 41300 73892
rect 41468 72548 41524 73836
rect 41244 71138 41300 71148
rect 41356 72492 41468 72548
rect 41132 70926 41134 70978
rect 41186 70926 41188 70978
rect 41132 70914 41188 70926
rect 41020 70756 41076 70766
rect 41356 70756 41412 72492
rect 41468 72482 41524 72492
rect 41580 73892 41748 73948
rect 41804 73948 41860 76974
rect 41916 75236 41972 79200
rect 42588 77138 42644 79200
rect 42588 77086 42590 77138
rect 42642 77086 42644 77138
rect 42588 77074 42644 77086
rect 42700 77026 42756 77038
rect 42700 76974 42702 77026
rect 42754 76974 42756 77026
rect 42700 76578 42756 76974
rect 42700 76526 42702 76578
rect 42754 76526 42756 76578
rect 42700 76514 42756 76526
rect 43260 76580 43316 79200
rect 43708 77364 43764 77374
rect 43260 76524 43428 76580
rect 42812 76356 42868 76366
rect 41916 75170 41972 75180
rect 42252 75570 42308 75582
rect 42252 75518 42254 75570
rect 42306 75518 42308 75570
rect 42252 74900 42308 75518
rect 42476 75460 42532 75470
rect 42700 75460 42756 75470
rect 42812 75460 42868 76300
rect 42476 75458 42644 75460
rect 42476 75406 42478 75458
rect 42530 75406 42644 75458
rect 42476 75404 42644 75406
rect 42476 75394 42532 75404
rect 42252 74834 42308 74844
rect 42476 75236 42532 75246
rect 42476 74898 42532 75180
rect 42476 74846 42478 74898
rect 42530 74846 42532 74898
rect 42028 74676 42084 74686
rect 42028 74226 42084 74620
rect 42028 74174 42030 74226
rect 42082 74174 42084 74226
rect 42028 74162 42084 74174
rect 42140 74116 42196 74126
rect 42140 74002 42196 74060
rect 42476 74116 42532 74846
rect 42476 74050 42532 74060
rect 42588 74898 42644 75404
rect 42700 75458 42868 75460
rect 42700 75406 42702 75458
rect 42754 75406 42868 75458
rect 42700 75404 42868 75406
rect 42700 75394 42756 75404
rect 42588 74846 42590 74898
rect 42642 74846 42644 74898
rect 42140 73950 42142 74002
rect 42194 73950 42196 74002
rect 41804 73892 42084 73948
rect 42140 73938 42196 73950
rect 42588 73948 42644 74846
rect 42700 74900 42756 74910
rect 42700 74806 42756 74844
rect 42812 74676 42868 75404
rect 42924 75570 42980 75582
rect 42924 75518 42926 75570
rect 42978 75518 42980 75570
rect 42924 75236 42980 75518
rect 43036 75572 43092 75582
rect 43036 75478 43092 75516
rect 43260 75572 43316 75582
rect 42924 75170 42980 75180
rect 43148 75124 43204 75134
rect 43148 75030 43204 75068
rect 41580 71202 41636 73892
rect 41692 73218 41748 73230
rect 41692 73166 41694 73218
rect 41746 73166 41748 73218
rect 41692 72660 41748 73166
rect 41692 72594 41748 72604
rect 41692 72324 41748 72334
rect 41692 72230 41748 72268
rect 41580 71150 41582 71202
rect 41634 71150 41636 71202
rect 41580 71138 41636 71150
rect 41804 71764 41860 71774
rect 41804 71092 41860 71708
rect 42028 71092 42084 73892
rect 42252 73892 42644 73948
rect 42700 74620 42868 74676
rect 43148 74788 43204 74798
rect 42252 73554 42308 73892
rect 42700 73780 42756 74620
rect 42924 74114 42980 74126
rect 42924 74062 42926 74114
rect 42978 74062 42980 74114
rect 42700 73714 42756 73724
rect 42812 74004 42868 74014
rect 42252 73502 42254 73554
rect 42306 73502 42308 73554
rect 42252 73490 42308 73502
rect 42700 73220 42756 73230
rect 42700 73126 42756 73164
rect 42812 72546 42868 73948
rect 42924 73780 42980 74062
rect 43148 74114 43204 74732
rect 43148 74062 43150 74114
rect 43202 74062 43204 74114
rect 43148 74050 43204 74062
rect 42924 73714 42980 73724
rect 43260 73444 43316 75516
rect 43372 73668 43428 76524
rect 43708 76468 43764 77308
rect 43820 76692 43876 76702
rect 43820 76598 43876 76636
rect 43708 76412 43876 76468
rect 43708 76242 43764 76254
rect 43708 76190 43710 76242
rect 43762 76190 43764 76242
rect 43708 75684 43764 76190
rect 43596 75628 43764 75684
rect 43484 75572 43540 75582
rect 43484 75478 43540 75516
rect 43596 75348 43652 75628
rect 43820 75570 43876 76412
rect 43932 75684 43988 79200
rect 44380 77138 44436 77150
rect 44380 77086 44382 77138
rect 44434 77086 44436 77138
rect 44044 76244 44100 76254
rect 44044 76150 44100 76188
rect 43932 75618 43988 75628
rect 43820 75518 43822 75570
rect 43874 75518 43876 75570
rect 43820 75506 43876 75518
rect 43708 75460 43764 75498
rect 43708 75394 43764 75404
rect 43932 75458 43988 75470
rect 43932 75406 43934 75458
rect 43986 75406 43988 75458
rect 43596 75282 43652 75292
rect 43708 75236 43764 75246
rect 43708 75012 43764 75180
rect 43932 75124 43988 75406
rect 43932 75058 43988 75068
rect 44044 75458 44100 75470
rect 44044 75406 44046 75458
rect 44098 75406 44100 75458
rect 43372 73602 43428 73612
rect 43484 75010 43764 75012
rect 43484 74958 43710 75010
rect 43762 74958 43764 75010
rect 43484 74956 43764 74958
rect 43484 74004 43540 74956
rect 43708 74946 43764 74956
rect 43932 74898 43988 74910
rect 43932 74846 43934 74898
rect 43986 74846 43988 74898
rect 43820 74788 43876 74798
rect 43820 74694 43876 74732
rect 43260 73388 43428 73444
rect 43148 73332 43204 73342
rect 43148 73238 43204 73276
rect 42924 73108 42980 73118
rect 42980 73052 43092 73108
rect 42924 72976 42980 73052
rect 42812 72494 42814 72546
rect 42866 72494 42868 72546
rect 42812 72482 42868 72494
rect 42252 72434 42308 72446
rect 42252 72382 42254 72434
rect 42306 72382 42308 72434
rect 42252 71652 42308 72382
rect 43036 71986 43092 73052
rect 43372 72996 43428 73388
rect 43036 71934 43038 71986
rect 43090 71934 43092 71986
rect 43036 71922 43092 71934
rect 43148 72660 43204 72670
rect 42924 71876 42980 71886
rect 42252 71586 42308 71596
rect 42812 71762 42868 71774
rect 42812 71710 42814 71762
rect 42866 71710 42868 71762
rect 42812 71652 42868 71710
rect 42812 71586 42868 71596
rect 42140 71092 42196 71102
rect 42028 71090 42196 71092
rect 42028 71038 42142 71090
rect 42194 71038 42196 71090
rect 42028 71036 42196 71038
rect 41804 71026 41860 71036
rect 42140 71026 42196 71036
rect 42812 70980 42868 70990
rect 42812 70886 42868 70924
rect 41076 70700 41412 70756
rect 41020 70418 41076 70700
rect 41020 70366 41022 70418
rect 41074 70366 41076 70418
rect 41020 70354 41076 70366
rect 42812 70420 42868 70430
rect 42924 70420 42980 71820
rect 42812 70418 42980 70420
rect 42812 70366 42814 70418
rect 42866 70366 42980 70418
rect 42812 70364 42980 70366
rect 42812 70354 42868 70364
rect 40460 70254 40462 70306
rect 40514 70254 40516 70306
rect 40460 70242 40516 70254
rect 39676 69470 39678 69522
rect 39730 69470 39732 69522
rect 39004 69458 39060 69468
rect 39676 69458 39732 69470
rect 40124 70196 40180 70206
rect 40124 69522 40180 70140
rect 43148 70194 43204 72604
rect 43260 71876 43316 71886
rect 43260 71782 43316 71820
rect 43372 71652 43428 72940
rect 43148 70142 43150 70194
rect 43202 70142 43204 70194
rect 43148 70130 43204 70142
rect 43260 71596 43428 71652
rect 40124 69470 40126 69522
rect 40178 69470 40180 69522
rect 40124 69458 40180 69470
rect 43260 69522 43316 71596
rect 43372 70196 43428 70206
rect 43484 70196 43540 73948
rect 43708 74676 43764 74686
rect 43596 72436 43652 72446
rect 43596 71762 43652 72380
rect 43596 71710 43598 71762
rect 43650 71710 43652 71762
rect 43596 71698 43652 71710
rect 43596 71428 43652 71438
rect 43596 70978 43652 71372
rect 43596 70926 43598 70978
rect 43650 70926 43652 70978
rect 43596 70914 43652 70926
rect 43372 70194 43540 70196
rect 43372 70142 43374 70194
rect 43426 70142 43540 70194
rect 43372 70140 43540 70142
rect 43372 70130 43428 70140
rect 43708 69970 43764 74620
rect 43932 74228 43988 74846
rect 44044 74340 44100 75406
rect 44156 75460 44212 75470
rect 44156 75012 44212 75404
rect 44156 74898 44212 74956
rect 44156 74846 44158 74898
rect 44210 74846 44212 74898
rect 44156 74834 44212 74846
rect 44268 75236 44324 75246
rect 44044 74274 44100 74284
rect 44268 74338 44324 75180
rect 44380 74676 44436 77086
rect 44604 76804 44660 79200
rect 44492 76748 44660 76804
rect 44828 77138 44884 77150
rect 44828 77086 44830 77138
rect 44882 77086 44884 77138
rect 44492 75572 44548 76748
rect 44492 75506 44548 75516
rect 44604 76578 44660 76590
rect 44604 76526 44606 76578
rect 44658 76526 44660 76578
rect 44604 75236 44660 76526
rect 44828 76466 44884 77086
rect 44828 76414 44830 76466
rect 44882 76414 44884 76466
rect 44828 76402 44884 76414
rect 45052 76580 45108 76590
rect 44604 75170 44660 75180
rect 44716 76244 44772 76254
rect 44716 75906 44772 76188
rect 44716 75854 44718 75906
rect 44770 75854 44772 75906
rect 44492 74900 44548 74910
rect 44492 74898 44660 74900
rect 44492 74846 44494 74898
rect 44546 74846 44660 74898
rect 44492 74844 44660 74846
rect 44492 74834 44548 74844
rect 44380 74610 44436 74620
rect 44604 74674 44660 74844
rect 44604 74622 44606 74674
rect 44658 74622 44660 74674
rect 44604 74610 44660 74622
rect 44268 74286 44270 74338
rect 44322 74286 44324 74338
rect 44268 74274 44324 74286
rect 44380 74452 44436 74462
rect 43932 74134 43988 74172
rect 44156 74116 44212 74154
rect 44156 74050 44212 74060
rect 44380 73948 44436 74396
rect 44716 73948 44772 75854
rect 45052 75908 45108 76524
rect 44828 75796 44884 75806
rect 44828 75702 44884 75740
rect 44940 75460 44996 75470
rect 44828 75458 44996 75460
rect 44828 75406 44942 75458
rect 44994 75406 44996 75458
rect 44828 75404 44996 75406
rect 44828 75236 44884 75404
rect 44940 75394 44996 75404
rect 44828 74564 44884 75180
rect 44940 75124 44996 75134
rect 45052 75124 45108 75852
rect 44940 75122 45108 75124
rect 44940 75070 44942 75122
rect 44994 75070 45108 75122
rect 44940 75068 45108 75070
rect 44940 75058 44996 75068
rect 45164 74788 45220 74798
rect 44828 74498 44884 74508
rect 44940 74674 44996 74686
rect 44940 74622 44942 74674
rect 44994 74622 44996 74674
rect 44828 74228 44884 74238
rect 44828 74134 44884 74172
rect 43820 73892 43876 73902
rect 43820 70420 43876 73836
rect 44156 73892 44212 73902
rect 44044 73556 44100 73566
rect 43932 73332 43988 73342
rect 43932 72658 43988 73276
rect 43932 72606 43934 72658
rect 43986 72606 43988 72658
rect 43932 72594 43988 72606
rect 43932 72436 43988 72446
rect 44044 72436 44100 73500
rect 44156 73330 44212 73836
rect 44268 73890 44324 73902
rect 44380 73892 44548 73948
rect 44716 73892 44884 73948
rect 44268 73838 44270 73890
rect 44322 73838 44324 73890
rect 44268 73780 44324 73838
rect 44268 73714 44324 73724
rect 44156 73278 44158 73330
rect 44210 73278 44212 73330
rect 44156 72772 44212 73278
rect 44380 73332 44436 73342
rect 44492 73332 44548 73892
rect 44716 73780 44772 73790
rect 44604 73444 44660 73454
rect 44604 73350 44660 73388
rect 44716 73442 44772 73724
rect 44716 73390 44718 73442
rect 44770 73390 44772 73442
rect 44716 73378 44772 73390
rect 44380 73330 44548 73332
rect 44380 73278 44382 73330
rect 44434 73278 44548 73330
rect 44380 73276 44548 73278
rect 44380 73266 44436 73276
rect 44156 72706 44212 72716
rect 43988 72380 44100 72436
rect 44156 72436 44212 72446
rect 44716 72436 44772 72446
rect 44156 72434 44772 72436
rect 44156 72382 44158 72434
rect 44210 72382 44718 72434
rect 44770 72382 44772 72434
rect 44156 72380 44772 72382
rect 43932 72304 43988 72380
rect 43932 71876 43988 71886
rect 44156 71876 44212 72380
rect 44716 72370 44772 72380
rect 43932 71874 44212 71876
rect 43932 71822 43934 71874
rect 43986 71822 44212 71874
rect 43932 71820 44212 71822
rect 43932 70980 43988 71820
rect 44492 71764 44548 71774
rect 44492 71670 44548 71708
rect 44716 71650 44772 71662
rect 44716 71598 44718 71650
rect 44770 71598 44772 71650
rect 44716 71428 44772 71598
rect 44716 71362 44772 71372
rect 44828 71204 44884 73892
rect 44940 73780 44996 74622
rect 44940 73714 44996 73724
rect 44940 73108 44996 73118
rect 44940 73014 44996 73052
rect 45164 72772 45220 74732
rect 45276 73948 45332 79200
rect 45836 77476 45892 77486
rect 45500 76580 45556 76590
rect 45500 76486 45556 76524
rect 45836 76578 45892 77420
rect 45836 76526 45838 76578
rect 45890 76526 45892 76578
rect 45836 76514 45892 76526
rect 45948 76468 46004 79200
rect 46620 77026 46676 79200
rect 46956 77476 47012 77486
rect 46620 76974 46622 77026
rect 46674 76974 46676 77026
rect 46620 76962 46676 76974
rect 46844 77026 46900 77038
rect 46844 76974 46846 77026
rect 46898 76974 46900 77026
rect 45948 76402 46004 76412
rect 46396 76356 46452 76366
rect 46396 76262 46452 76300
rect 46732 76242 46788 76254
rect 46732 76190 46734 76242
rect 46786 76190 46788 76242
rect 45500 76020 45556 76030
rect 45500 74676 45556 75964
rect 46732 75684 46788 76190
rect 46060 75682 46788 75684
rect 46060 75630 46734 75682
rect 46786 75630 46788 75682
rect 46060 75628 46788 75630
rect 45948 75570 46004 75582
rect 45948 75518 45950 75570
rect 46002 75518 46004 75570
rect 45612 75460 45668 75470
rect 45612 75366 45668 75404
rect 45948 75460 46004 75518
rect 45948 75394 46004 75404
rect 45948 75124 46004 75134
rect 46060 75124 46116 75628
rect 46732 75618 46788 75628
rect 46508 75458 46564 75470
rect 46844 75460 46900 76974
rect 46956 76692 47012 77420
rect 46956 76636 47124 76692
rect 46508 75406 46510 75458
rect 46562 75406 46564 75458
rect 46508 75236 46564 75406
rect 46508 75170 46564 75180
rect 46732 75404 46900 75460
rect 46956 76468 47012 76478
rect 45948 75122 46116 75124
rect 45948 75070 45950 75122
rect 46002 75070 46116 75122
rect 45948 75068 46116 75070
rect 45948 75058 46004 75068
rect 45724 74900 45780 74910
rect 45724 74806 45780 74844
rect 45500 74114 45556 74620
rect 45500 74062 45502 74114
rect 45554 74062 45556 74114
rect 45500 74050 45556 74062
rect 45836 74786 45892 74798
rect 45836 74734 45838 74786
rect 45890 74734 45892 74786
rect 45612 74004 45668 74042
rect 45276 73892 45444 73948
rect 45612 73938 45668 73948
rect 45724 74002 45780 74014
rect 45724 73950 45726 74002
rect 45778 73950 45780 74002
rect 45164 72716 45332 72772
rect 45164 72548 45220 72558
rect 45164 72454 45220 72492
rect 45052 72436 45108 72446
rect 44940 71762 44996 71774
rect 44940 71710 44942 71762
rect 44994 71710 44996 71762
rect 44940 71540 44996 71710
rect 44940 71474 44996 71484
rect 44380 71148 44884 71204
rect 44268 70980 44324 70990
rect 43932 70978 44324 70980
rect 43932 70926 44270 70978
rect 44322 70926 44324 70978
rect 43932 70924 44324 70926
rect 44268 70914 44324 70924
rect 43932 70420 43988 70430
rect 43820 70418 43988 70420
rect 43820 70366 43934 70418
rect 43986 70366 43988 70418
rect 43820 70364 43988 70366
rect 43932 70354 43988 70364
rect 44268 70420 44324 70430
rect 44380 70420 44436 71148
rect 45052 71092 45108 72380
rect 45164 71876 45220 71886
rect 45164 71782 45220 71820
rect 45276 71652 45332 72716
rect 45388 71988 45444 73892
rect 45724 73556 45780 73950
rect 45724 73490 45780 73500
rect 45612 73444 45668 73454
rect 45500 73218 45556 73230
rect 45500 73166 45502 73218
rect 45554 73166 45556 73218
rect 45500 72660 45556 73166
rect 45500 72594 45556 72604
rect 45612 72658 45668 73388
rect 45836 73218 45892 74734
rect 46060 74114 46116 75068
rect 46284 74900 46340 74910
rect 46060 74062 46062 74114
rect 46114 74062 46116 74114
rect 46060 74050 46116 74062
rect 46172 74786 46228 74798
rect 46172 74734 46174 74786
rect 46226 74734 46228 74786
rect 45836 73166 45838 73218
rect 45890 73166 45892 73218
rect 45836 73154 45892 73166
rect 45948 73780 46004 73790
rect 45948 73330 46004 73724
rect 46172 73556 46228 74734
rect 46172 73490 46228 73500
rect 46284 73892 46340 74844
rect 46396 74676 46452 74686
rect 46452 74620 46564 74676
rect 46396 74582 46452 74620
rect 45948 73278 45950 73330
rect 46002 73278 46004 73330
rect 45612 72606 45614 72658
rect 45666 72606 45668 72658
rect 45612 72594 45668 72606
rect 45724 71988 45780 71998
rect 45388 71986 45780 71988
rect 45388 71934 45726 71986
rect 45778 71934 45780 71986
rect 45388 71932 45780 71934
rect 45724 71922 45780 71932
rect 45948 71762 46004 73278
rect 45948 71710 45950 71762
rect 46002 71710 46004 71762
rect 45948 71698 46004 71710
rect 46060 73332 46116 73342
rect 44268 70418 44436 70420
rect 44268 70366 44270 70418
rect 44322 70366 44436 70418
rect 44268 70364 44436 70366
rect 44268 70354 44324 70364
rect 43708 69918 43710 69970
rect 43762 69918 43764 69970
rect 43708 69906 43764 69918
rect 43260 69470 43262 69522
rect 43314 69470 43316 69522
rect 43260 69458 43316 69470
rect 44380 69524 44436 70364
rect 44828 70980 44884 70990
rect 44828 70418 44884 70924
rect 44940 70980 44996 70990
rect 45052 70980 45108 71036
rect 44940 70978 45108 70980
rect 44940 70926 44942 70978
rect 44994 70926 45108 70978
rect 44940 70924 45108 70926
rect 45164 71596 45332 71652
rect 44940 70914 44996 70924
rect 45164 70532 45220 71596
rect 46060 71540 46116 73276
rect 46284 73332 46340 73836
rect 46284 73266 46340 73276
rect 46284 73108 46340 73118
rect 46284 72546 46340 73052
rect 46284 72494 46286 72546
rect 46338 72494 46340 72546
rect 46284 72482 46340 72494
rect 46396 72436 46452 72446
rect 46284 72324 46340 72334
rect 45724 71538 46116 71540
rect 45724 71486 46062 71538
rect 46114 71486 46116 71538
rect 45724 71484 46116 71486
rect 45612 71202 45668 71214
rect 45612 71150 45614 71202
rect 45666 71150 45668 71202
rect 45612 71092 45668 71150
rect 45612 70998 45668 71036
rect 45276 70532 45332 70542
rect 45164 70476 45276 70532
rect 44828 70366 44830 70418
rect 44882 70366 44884 70418
rect 44828 70354 44884 70366
rect 45276 70418 45332 70476
rect 45276 70366 45278 70418
rect 45330 70366 45332 70418
rect 45276 70354 45332 70366
rect 45724 70418 45780 71484
rect 46060 71474 46116 71484
rect 46172 71762 46228 71774
rect 46172 71710 46174 71762
rect 46226 71710 46228 71762
rect 46060 71204 46116 71214
rect 46060 71090 46116 71148
rect 46060 71038 46062 71090
rect 46114 71038 46116 71090
rect 46060 71026 46116 71038
rect 46172 70980 46228 71710
rect 46284 71650 46340 72268
rect 46284 71598 46286 71650
rect 46338 71598 46340 71650
rect 46284 71202 46340 71598
rect 46284 71150 46286 71202
rect 46338 71150 46340 71202
rect 46284 71138 46340 71150
rect 46396 71204 46452 72380
rect 46508 71988 46564 74620
rect 46620 73890 46676 73902
rect 46620 73838 46622 73890
rect 46674 73838 46676 73890
rect 46620 73668 46676 73838
rect 46620 73602 46676 73612
rect 46620 72548 46676 72558
rect 46620 72454 46676 72492
rect 46732 71988 46788 75404
rect 46844 74898 46900 74910
rect 46844 74846 46846 74898
rect 46898 74846 46900 74898
rect 46844 73108 46900 74846
rect 46844 73042 46900 73052
rect 46956 72436 47012 76412
rect 47068 75122 47124 76636
rect 47068 75070 47070 75122
rect 47122 75070 47124 75122
rect 47068 74004 47124 75070
rect 47180 75460 47236 75470
rect 47180 75010 47236 75404
rect 47180 74958 47182 75010
rect 47234 74958 47236 75010
rect 47180 74946 47236 74958
rect 47292 74116 47348 79200
rect 47404 75572 47460 75582
rect 47460 75516 47572 75572
rect 47404 75478 47460 75516
rect 47292 74050 47348 74060
rect 47404 75348 47460 75358
rect 47068 73938 47124 73948
rect 47292 73892 47348 73902
rect 47404 73892 47460 75292
rect 47292 73890 47460 73892
rect 47292 73838 47294 73890
rect 47346 73838 47460 73890
rect 47292 73836 47460 73838
rect 47292 73826 47348 73836
rect 47180 73444 47236 73454
rect 47180 73350 47236 73388
rect 47068 73332 47124 73342
rect 47068 72660 47124 73276
rect 47292 73330 47348 73342
rect 47292 73278 47294 73330
rect 47346 73278 47348 73330
rect 47180 73220 47236 73230
rect 47180 73106 47236 73164
rect 47180 73054 47182 73106
rect 47234 73054 47236 73106
rect 47180 73042 47236 73054
rect 47068 72604 47236 72660
rect 47068 72436 47124 72446
rect 46956 72434 47124 72436
rect 46956 72382 47070 72434
rect 47122 72382 47124 72434
rect 46956 72380 47124 72382
rect 47068 72370 47124 72380
rect 46508 71922 46564 71932
rect 46620 71932 46788 71988
rect 47180 71988 47236 72604
rect 47292 72548 47348 73278
rect 47292 72482 47348 72492
rect 47180 71986 47460 71988
rect 47180 71934 47182 71986
rect 47234 71934 47460 71986
rect 47180 71932 47460 71934
rect 46396 71138 46452 71148
rect 46508 71202 46564 71214
rect 46508 71150 46510 71202
rect 46562 71150 46564 71202
rect 46508 70980 46564 71150
rect 46228 70978 46564 70980
rect 46228 70926 46510 70978
rect 46562 70926 46564 70978
rect 46228 70924 46564 70926
rect 46172 70848 46228 70924
rect 46508 70914 46564 70924
rect 45724 70366 45726 70418
rect 45778 70366 45780 70418
rect 45724 70354 45780 70366
rect 46172 70420 46228 70430
rect 46172 70326 46228 70364
rect 46620 70418 46676 71932
rect 47180 71922 47236 71932
rect 46732 71650 46788 71662
rect 46732 71598 46734 71650
rect 46786 71598 46788 71650
rect 46732 71538 46788 71598
rect 46732 71486 46734 71538
rect 46786 71486 46788 71538
rect 46732 71474 46788 71486
rect 46956 71202 47012 71214
rect 46956 71150 46958 71202
rect 47010 71150 47012 71202
rect 46956 71090 47012 71150
rect 46956 71038 46958 71090
rect 47010 71038 47012 71090
rect 46956 71026 47012 71038
rect 47404 71090 47460 71932
rect 47404 71038 47406 71090
rect 47458 71038 47460 71090
rect 47404 71026 47460 71038
rect 46620 70366 46622 70418
rect 46674 70366 46676 70418
rect 46620 70354 46676 70366
rect 47180 70420 47236 70430
rect 47516 70420 47572 75516
rect 47740 75460 47796 75470
rect 47628 75458 47796 75460
rect 47628 75406 47742 75458
rect 47794 75406 47796 75458
rect 47628 75404 47796 75406
rect 47628 72324 47684 75404
rect 47740 75394 47796 75404
rect 47852 74228 47908 74266
rect 47852 74162 47908 74172
rect 47852 74004 47908 74014
rect 47852 73780 47908 73948
rect 47964 73948 48020 79200
rect 48524 76580 48580 76590
rect 48412 76020 48468 76030
rect 48412 75794 48468 75964
rect 48412 75742 48414 75794
rect 48466 75742 48468 75794
rect 48412 75730 48468 75742
rect 48300 75460 48356 75470
rect 48300 75366 48356 75404
rect 48524 75236 48580 76524
rect 48412 75180 48580 75236
rect 48188 74676 48244 74686
rect 48188 74674 48356 74676
rect 48188 74622 48190 74674
rect 48242 74622 48356 74674
rect 48188 74620 48356 74622
rect 48188 74610 48244 74620
rect 47964 73892 48244 73948
rect 47852 73724 48020 73780
rect 47852 73556 47908 73566
rect 47852 73462 47908 73500
rect 47964 73218 48020 73724
rect 47964 73166 47966 73218
rect 48018 73166 48020 73218
rect 47628 72230 47684 72268
rect 47740 72548 47796 72558
rect 47628 71988 47684 71998
rect 47740 71988 47796 72492
rect 47628 71986 47796 71988
rect 47628 71934 47630 71986
rect 47682 71934 47796 71986
rect 47628 71932 47796 71934
rect 47852 71988 47908 71998
rect 47628 71922 47684 71932
rect 47852 71092 47908 71932
rect 47964 71538 48020 73166
rect 48188 72434 48244 73892
rect 48188 72382 48190 72434
rect 48242 72382 48244 72434
rect 48188 72370 48244 72382
rect 48300 72324 48356 74620
rect 48412 72548 48468 75180
rect 48636 75012 48692 79200
rect 48860 77026 48916 77038
rect 48860 76974 48862 77026
rect 48914 76974 48916 77026
rect 48860 76578 48916 76974
rect 48860 76526 48862 76578
rect 48914 76526 48916 76578
rect 48860 76514 48916 76526
rect 49084 76356 49140 76366
rect 48972 76132 49028 76142
rect 48972 75794 49028 76076
rect 48972 75742 48974 75794
rect 49026 75742 49028 75794
rect 48972 75730 49028 75742
rect 49084 75796 49140 76300
rect 49084 75682 49140 75740
rect 49084 75630 49086 75682
rect 49138 75630 49140 75682
rect 49084 75618 49140 75630
rect 49084 75460 49140 75470
rect 48636 74946 48692 74956
rect 48748 75124 48804 75134
rect 48524 74674 48580 74686
rect 48524 74622 48526 74674
rect 48578 74622 48580 74674
rect 48524 74340 48580 74622
rect 48636 74340 48692 74350
rect 48524 74338 48692 74340
rect 48524 74286 48638 74338
rect 48690 74286 48692 74338
rect 48524 74284 48692 74286
rect 48636 74274 48692 74284
rect 48524 74116 48580 74126
rect 48524 73554 48580 74060
rect 48748 74114 48804 75068
rect 48748 74062 48750 74114
rect 48802 74062 48804 74114
rect 48748 74050 48804 74062
rect 48860 75010 48916 75022
rect 49084 75012 49140 75404
rect 48860 74958 48862 75010
rect 48914 74958 48916 75010
rect 48636 73892 48692 73902
rect 48636 73798 48692 73836
rect 48524 73502 48526 73554
rect 48578 73502 48580 73554
rect 48524 73490 48580 73502
rect 48860 73444 48916 74958
rect 48860 73378 48916 73388
rect 48972 75010 49140 75012
rect 48972 74958 49086 75010
rect 49138 74958 49140 75010
rect 48972 74956 49140 74958
rect 48412 72482 48468 72492
rect 48300 72268 48468 72324
rect 48076 71988 48132 71998
rect 48076 71894 48132 71932
rect 47964 71486 47966 71538
rect 48018 71486 48020 71538
rect 47964 71474 48020 71486
rect 48412 71316 48468 72268
rect 48972 71876 49028 74956
rect 49084 74946 49140 74956
rect 49308 74900 49364 79200
rect 49980 76692 50036 79200
rect 50652 77028 50708 79200
rect 50652 76962 50708 76972
rect 50556 76860 50820 76870
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50556 76794 50820 76804
rect 49980 76636 50260 76692
rect 49868 76578 49924 76590
rect 49868 76526 49870 76578
rect 49922 76526 49924 76578
rect 49756 76244 49812 76254
rect 49420 76242 49812 76244
rect 49420 76190 49758 76242
rect 49810 76190 49812 76242
rect 49420 76188 49812 76190
rect 49420 75570 49476 76188
rect 49756 76178 49812 76188
rect 49868 75684 49924 76526
rect 49420 75518 49422 75570
rect 49474 75518 49476 75570
rect 49420 75506 49476 75518
rect 49532 75628 49924 75684
rect 50092 76466 50148 76478
rect 50092 76414 50094 76466
rect 50146 76414 50148 76466
rect 49532 75458 49588 75628
rect 49532 75406 49534 75458
rect 49586 75406 49588 75458
rect 49532 75348 49588 75406
rect 49756 75460 49812 75470
rect 49756 75366 49812 75404
rect 49196 74844 49364 74900
rect 49420 75292 49588 75348
rect 49196 73948 49252 74844
rect 49308 74340 49364 74350
rect 49308 74246 49364 74284
rect 49084 73892 49252 73948
rect 49084 72434 49140 73892
rect 49420 73444 49476 75292
rect 49420 73378 49476 73388
rect 49532 75012 49588 75022
rect 49980 75012 50036 75022
rect 49420 73220 49476 73230
rect 49420 73126 49476 73164
rect 49084 72382 49086 72434
rect 49138 72382 49140 72434
rect 49084 72370 49140 72382
rect 49420 71876 49476 71886
rect 48972 71874 49476 71876
rect 48972 71822 49422 71874
rect 49474 71822 49476 71874
rect 48972 71820 49476 71822
rect 49420 71810 49476 71820
rect 48412 71250 48468 71260
rect 48524 71650 48580 71662
rect 48524 71598 48526 71650
rect 48578 71598 48580 71650
rect 48524 71538 48580 71598
rect 48524 71486 48526 71538
rect 48578 71486 48580 71538
rect 47852 70960 47908 71036
rect 47180 70418 47572 70420
rect 47180 70366 47182 70418
rect 47234 70366 47572 70418
rect 47180 70364 47572 70366
rect 48300 70756 48356 70766
rect 48524 70756 48580 71486
rect 48748 71092 48804 71102
rect 48748 70998 48804 71036
rect 49308 71092 49364 71102
rect 49308 70998 49364 71036
rect 48300 70754 48580 70756
rect 48300 70702 48302 70754
rect 48354 70702 48580 70754
rect 48300 70700 48580 70702
rect 48300 70420 48356 70700
rect 49532 70420 49588 74956
rect 49644 75010 50036 75012
rect 49644 74958 49982 75010
rect 50034 74958 50036 75010
rect 49644 74956 50036 74958
rect 49644 73332 49700 74956
rect 49980 74946 50036 74956
rect 50092 74788 50148 76414
rect 49980 74732 50148 74788
rect 49644 73266 49700 73276
rect 49756 74116 49812 74126
rect 49756 74002 49812 74060
rect 49756 73950 49758 74002
rect 49810 73950 49812 74002
rect 49644 73106 49700 73118
rect 49644 73054 49646 73106
rect 49698 73054 49700 73106
rect 49644 72660 49700 73054
rect 49644 72546 49700 72604
rect 49756 72658 49812 73950
rect 49868 74004 49924 74042
rect 49868 73938 49924 73948
rect 49980 73892 50036 74732
rect 50092 74228 50148 74238
rect 50092 74114 50148 74172
rect 50092 74062 50094 74114
rect 50146 74062 50148 74114
rect 50092 74050 50148 74062
rect 49980 73826 50036 73836
rect 49868 73108 49924 73118
rect 49868 73106 50148 73108
rect 49868 73054 49870 73106
rect 49922 73054 50148 73106
rect 49868 73052 50148 73054
rect 49868 73042 49924 73052
rect 49756 72606 49758 72658
rect 49810 72606 49812 72658
rect 49756 72594 49812 72606
rect 49868 72884 49924 72894
rect 49644 72494 49646 72546
rect 49698 72494 49700 72546
rect 49644 72482 49700 72494
rect 49868 72546 49924 72828
rect 49868 72494 49870 72546
rect 49922 72494 49924 72546
rect 49868 72482 49924 72494
rect 50092 72548 50148 73052
rect 50092 72434 50148 72492
rect 50092 72382 50094 72434
rect 50146 72382 50148 72434
rect 50092 72370 50148 72382
rect 49868 72324 49924 72334
rect 49644 70754 49700 70766
rect 49644 70702 49646 70754
rect 49698 70702 49700 70754
rect 49644 70644 49700 70702
rect 49868 70644 49924 72268
rect 50204 71988 50260 76636
rect 50316 76466 50372 76478
rect 50316 76414 50318 76466
rect 50370 76414 50372 76466
rect 50316 75124 50372 76414
rect 51100 76356 51156 76366
rect 51100 76354 51268 76356
rect 51100 76302 51102 76354
rect 51154 76302 51268 76354
rect 51100 76300 51268 76302
rect 51100 76290 51156 76300
rect 50316 75058 50372 75068
rect 50428 75682 50484 75694
rect 50428 75630 50430 75682
rect 50482 75630 50484 75682
rect 50316 74900 50372 74910
rect 50316 74806 50372 74844
rect 50316 74004 50372 74014
rect 50316 73554 50372 73948
rect 50316 73502 50318 73554
rect 50370 73502 50372 73554
rect 50316 73490 50372 73502
rect 50428 73444 50484 75630
rect 50876 75458 50932 75470
rect 50876 75406 50878 75458
rect 50930 75406 50932 75458
rect 50556 75292 50820 75302
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50556 75226 50820 75236
rect 50764 75012 50820 75022
rect 50764 74338 50820 74956
rect 50876 74900 50932 75406
rect 50988 75458 51044 75470
rect 50988 75406 50990 75458
rect 51042 75406 51044 75458
rect 50988 75124 51044 75406
rect 50988 75058 51044 75068
rect 51100 75458 51156 75470
rect 51100 75406 51102 75458
rect 51154 75406 51156 75458
rect 50876 74834 50932 74844
rect 50764 74286 50766 74338
rect 50818 74286 50820 74338
rect 50764 74274 50820 74286
rect 50988 74786 51044 74798
rect 50988 74734 50990 74786
rect 51042 74734 51044 74786
rect 50652 74116 50708 74126
rect 50652 74022 50708 74060
rect 50876 74004 50932 74042
rect 50876 73938 50932 73948
rect 50556 73724 50820 73734
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50556 73658 50820 73668
rect 50988 73556 51044 74734
rect 51100 74340 51156 75406
rect 51100 74274 51156 74284
rect 51212 74116 51268 76300
rect 51324 74676 51380 79200
rect 51548 77028 51604 77038
rect 51436 74900 51492 74910
rect 51436 74806 51492 74844
rect 51548 74788 51604 76972
rect 51996 76468 52052 79200
rect 51996 76402 52052 76412
rect 52668 76356 52724 79200
rect 53228 77252 53284 77262
rect 52892 77028 52948 77038
rect 52892 76578 52948 76972
rect 52892 76526 52894 76578
rect 52946 76526 52948 76578
rect 52892 76514 52948 76526
rect 52668 76290 52724 76300
rect 52332 76020 52388 76030
rect 52332 75682 52388 75964
rect 53116 75908 53172 75918
rect 53116 75814 53172 75852
rect 52332 75630 52334 75682
rect 52386 75630 52388 75682
rect 52332 75618 52388 75630
rect 53004 75684 53060 75694
rect 53004 75590 53060 75628
rect 51660 75458 51716 75470
rect 51660 75406 51662 75458
rect 51714 75406 51716 75458
rect 51660 75236 51716 75406
rect 51660 75170 51716 75180
rect 51772 75458 51828 75470
rect 51772 75406 51774 75458
rect 51826 75406 51828 75458
rect 51772 75012 51828 75406
rect 51884 75460 51940 75470
rect 51884 75458 52052 75460
rect 51884 75406 51886 75458
rect 51938 75406 52052 75458
rect 51884 75404 52052 75406
rect 51884 75394 51940 75404
rect 51548 74722 51604 74732
rect 51660 74956 51828 75012
rect 51324 74620 51492 74676
rect 51436 74564 51492 74620
rect 51436 74508 51604 74564
rect 51212 74050 51268 74060
rect 51324 74228 51380 74238
rect 51324 74114 51380 74172
rect 51324 74062 51326 74114
rect 51378 74062 51380 74114
rect 51324 74050 51380 74062
rect 51436 74116 51492 74126
rect 51100 74004 51156 74042
rect 51436 73948 51492 74060
rect 51100 73938 51156 73948
rect 51212 73892 51492 73948
rect 51212 73556 51268 73892
rect 51548 73668 51604 74508
rect 51548 73602 51604 73612
rect 51660 73556 51716 74956
rect 51996 74900 52052 75404
rect 52892 75458 52948 75470
rect 52892 75406 52894 75458
rect 52946 75406 52948 75458
rect 52668 75012 52724 75022
rect 52668 75010 52836 75012
rect 52668 74958 52670 75010
rect 52722 74958 52836 75010
rect 52668 74956 52836 74958
rect 52668 74946 52724 74956
rect 51884 74786 51940 74798
rect 51884 74734 51886 74786
rect 51938 74734 51940 74786
rect 51884 74116 51940 74734
rect 51884 74050 51940 74060
rect 51996 74564 52052 74844
rect 51996 74002 52052 74508
rect 52108 74340 52164 74350
rect 52108 74114 52164 74284
rect 52108 74062 52110 74114
rect 52162 74062 52164 74114
rect 52108 74050 52164 74062
rect 52780 74228 52836 74956
rect 52892 74676 52948 75406
rect 53004 75012 53060 75022
rect 53004 74918 53060 74956
rect 52892 74610 52948 74620
rect 51996 73950 51998 74002
rect 52050 73950 52052 74002
rect 51772 73892 51828 73902
rect 51772 73798 51828 73836
rect 50988 73500 51156 73556
rect 51212 73500 51492 73556
rect 51660 73500 51828 73556
rect 50876 73444 50932 73454
rect 50428 73442 50932 73444
rect 50428 73390 50878 73442
rect 50930 73390 50932 73442
rect 50428 73388 50932 73390
rect 50316 73332 50372 73342
rect 50876 73332 50932 73388
rect 51100 73442 51156 73500
rect 51100 73390 51102 73442
rect 51154 73390 51156 73442
rect 51100 73332 51156 73390
rect 51212 73332 51268 73342
rect 50876 73276 51044 73332
rect 51100 73330 51268 73332
rect 51100 73278 51214 73330
rect 51266 73278 51268 73330
rect 51100 73276 51268 73278
rect 50316 72324 50372 73276
rect 50764 73220 50820 73230
rect 50764 73126 50820 73164
rect 50876 72772 50932 72782
rect 50876 72658 50932 72716
rect 50876 72606 50878 72658
rect 50930 72606 50932 72658
rect 50876 72594 50932 72606
rect 50764 72548 50820 72558
rect 50764 72454 50820 72492
rect 50316 72258 50372 72268
rect 50988 72324 51044 73276
rect 51212 73266 51268 73276
rect 50988 72258 51044 72268
rect 51100 73108 51156 73118
rect 50556 72156 50820 72166
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50556 72090 50820 72100
rect 50204 71932 50372 71988
rect 50204 71764 50260 71774
rect 50204 71670 50260 71708
rect 50204 70868 50260 70878
rect 50316 70868 50372 71932
rect 50876 71092 50932 71102
rect 51100 71092 51156 73052
rect 51436 71876 51492 73500
rect 51548 73332 51604 73342
rect 51548 73330 51716 73332
rect 51548 73278 51550 73330
rect 51602 73278 51716 73330
rect 51548 73276 51716 73278
rect 51548 73266 51604 73276
rect 51548 72660 51604 72670
rect 51548 72566 51604 72604
rect 51660 72434 51716 73276
rect 51772 72772 51828 73500
rect 51996 73444 52052 73950
rect 52780 74002 52836 74172
rect 53228 74226 53284 77196
rect 53340 76692 53396 79200
rect 54012 77364 54068 79200
rect 54012 77298 54068 77308
rect 53340 76626 53396 76636
rect 53900 76580 53956 76590
rect 54684 76580 54740 79200
rect 55020 76580 55076 76590
rect 54684 76578 55076 76580
rect 54684 76526 55022 76578
rect 55074 76526 55076 76578
rect 54684 76524 55076 76526
rect 53900 76486 53956 76524
rect 54236 76466 54292 76478
rect 54236 76414 54238 76466
rect 54290 76414 54292 76466
rect 54236 76356 54292 76414
rect 54236 76290 54292 76300
rect 54348 76020 54404 76030
rect 53228 74174 53230 74226
rect 53282 74174 53284 74226
rect 53228 74162 53284 74174
rect 53564 75796 53620 75806
rect 53564 75010 53620 75740
rect 54124 75684 54180 75694
rect 54124 75590 54180 75628
rect 53788 75572 53844 75582
rect 53788 75478 53844 75516
rect 53564 74958 53566 75010
rect 53618 74958 53620 75010
rect 52780 73950 52782 74002
rect 52834 73950 52836 74002
rect 52780 73938 52836 73950
rect 52892 74114 52948 74126
rect 52892 74062 52894 74114
rect 52946 74062 52948 74114
rect 51996 73378 52052 73388
rect 52332 73668 52388 73678
rect 52108 73220 52164 73230
rect 51772 72706 51828 72716
rect 51996 73218 52164 73220
rect 51996 73166 52110 73218
rect 52162 73166 52164 73218
rect 51996 73164 52164 73166
rect 51996 72660 52052 73164
rect 52108 73154 52164 73164
rect 51884 72548 51940 72558
rect 51884 72454 51940 72492
rect 51660 72382 51662 72434
rect 51714 72382 51716 72434
rect 50932 71036 51156 71092
rect 51212 71820 51492 71876
rect 51548 72324 51604 72334
rect 50876 70960 50932 71036
rect 50204 70866 50372 70868
rect 50204 70814 50206 70866
rect 50258 70814 50372 70866
rect 50204 70812 50372 70814
rect 50204 70802 50260 70812
rect 49644 70588 49924 70644
rect 49756 70420 49812 70430
rect 49532 70418 49812 70420
rect 49532 70366 49758 70418
rect 49810 70366 49812 70418
rect 49532 70364 49812 70366
rect 49868 70420 49924 70588
rect 50556 70588 50820 70598
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50556 70522 50820 70532
rect 50204 70420 50260 70430
rect 49868 70364 50204 70420
rect 47180 70354 47236 70364
rect 48300 70354 48356 70364
rect 49756 70354 49812 70364
rect 50204 70288 50260 70364
rect 50652 70420 50708 70430
rect 50652 70326 50708 70364
rect 51100 70420 51156 70430
rect 51212 70420 51268 71820
rect 51548 71764 51604 72268
rect 51324 71762 51604 71764
rect 51324 71710 51550 71762
rect 51602 71710 51604 71762
rect 51324 71708 51604 71710
rect 51324 71090 51380 71708
rect 51548 71698 51604 71708
rect 51660 71650 51716 72382
rect 51996 72324 52052 72604
rect 51660 71598 51662 71650
rect 51714 71598 51716 71650
rect 51660 71586 51716 71598
rect 51772 72268 52052 72324
rect 52108 72548 52164 72558
rect 51324 71038 51326 71090
rect 51378 71038 51380 71090
rect 51324 71026 51380 71038
rect 51772 70978 51828 72268
rect 51884 71764 51940 71774
rect 51884 71090 51940 71708
rect 51884 71038 51886 71090
rect 51938 71038 51940 71090
rect 51884 71026 51940 71038
rect 51772 70926 51774 70978
rect 51826 70926 51828 70978
rect 51772 70914 51828 70926
rect 52108 70978 52164 72492
rect 52332 71986 52388 73612
rect 52892 73442 52948 74062
rect 52892 73390 52894 73442
rect 52946 73390 52948 73442
rect 52892 73378 52948 73390
rect 53116 73444 53172 73454
rect 52444 73330 52500 73342
rect 52444 73278 52446 73330
rect 52498 73278 52500 73330
rect 52444 72548 52500 73278
rect 52444 72416 52500 72492
rect 53004 72548 53060 72558
rect 52668 72436 52724 72446
rect 52332 71934 52334 71986
rect 52386 71934 52388 71986
rect 52332 71922 52388 71934
rect 52556 72380 52668 72436
rect 52556 71652 52612 72380
rect 52668 72342 52724 72380
rect 52108 70926 52110 70978
rect 52162 70926 52164 70978
rect 52108 70914 52164 70926
rect 52332 71596 52612 71652
rect 52892 72324 52948 72334
rect 52332 70978 52388 71596
rect 52892 71090 52948 72268
rect 53004 71874 53060 72492
rect 53004 71822 53006 71874
rect 53058 71822 53060 71874
rect 53004 71810 53060 71822
rect 52892 71038 52894 71090
rect 52946 71038 52948 71090
rect 52892 71026 52948 71038
rect 53116 71092 53172 73388
rect 53564 73330 53620 74958
rect 53900 75458 53956 75470
rect 53900 75406 53902 75458
rect 53954 75406 53956 75458
rect 53788 74898 53844 74910
rect 53788 74846 53790 74898
rect 53842 74846 53844 74898
rect 53788 74340 53844 74846
rect 53900 74340 53956 75406
rect 54012 75460 54068 75470
rect 54012 75012 54068 75404
rect 54348 75348 54404 75964
rect 54460 75684 54516 75694
rect 54460 75590 54516 75628
rect 54348 75292 54516 75348
rect 54348 75124 54404 75134
rect 54012 74898 54068 74956
rect 54012 74846 54014 74898
rect 54066 74846 54068 74898
rect 54012 74834 54068 74846
rect 54236 75122 54404 75124
rect 54236 75070 54350 75122
rect 54402 75070 54404 75122
rect 54236 75068 54404 75070
rect 53900 74284 54180 74340
rect 53564 73278 53566 73330
rect 53618 73278 53620 73330
rect 53564 72772 53620 73278
rect 53676 74228 53732 74238
rect 53676 73330 53732 74172
rect 53676 73278 53678 73330
rect 53730 73278 53732 73330
rect 53676 73266 53732 73278
rect 53788 73332 53844 74284
rect 53900 74116 53956 74126
rect 53900 74114 54068 74116
rect 53900 74062 53902 74114
rect 53954 74062 54068 74114
rect 53900 74060 54068 74062
rect 53900 74050 53956 74060
rect 54012 73442 54068 74060
rect 54124 73948 54180 74284
rect 54236 74114 54292 75068
rect 54348 75058 54404 75068
rect 54348 74900 54404 74910
rect 54348 74806 54404 74844
rect 54236 74062 54238 74114
rect 54290 74062 54292 74114
rect 54236 74050 54292 74062
rect 54124 73892 54292 73948
rect 54012 73390 54014 73442
rect 54066 73390 54068 73442
rect 54012 73378 54068 73390
rect 54124 73556 54180 73566
rect 53900 73332 53956 73342
rect 53788 73330 53956 73332
rect 53788 73278 53902 73330
rect 53954 73278 53956 73330
rect 53788 73276 53956 73278
rect 53900 73266 53956 73276
rect 53340 72660 53396 72670
rect 53228 72548 53284 72558
rect 53228 71762 53284 72492
rect 53340 72546 53396 72604
rect 53340 72494 53342 72546
rect 53394 72494 53396 72546
rect 53340 72482 53396 72494
rect 53228 71710 53230 71762
rect 53282 71710 53284 71762
rect 53228 71698 53284 71710
rect 53564 71762 53620 72716
rect 53564 71710 53566 71762
rect 53618 71710 53620 71762
rect 53564 71698 53620 71710
rect 54124 72324 54180 73500
rect 53228 71092 53284 71102
rect 53116 71090 53284 71092
rect 53116 71038 53230 71090
rect 53282 71038 53284 71090
rect 53116 71036 53284 71038
rect 52332 70926 52334 70978
rect 52386 70926 52388 70978
rect 52332 70914 52388 70926
rect 52556 70532 52612 70542
rect 51100 70418 51268 70420
rect 51100 70366 51102 70418
rect 51154 70366 51268 70418
rect 51100 70364 51268 70366
rect 51660 70420 51716 70430
rect 51100 70354 51156 70364
rect 51660 70326 51716 70364
rect 52556 70418 52612 70476
rect 52556 70366 52558 70418
rect 52610 70366 52612 70418
rect 52556 70354 52612 70366
rect 53004 70420 53060 70430
rect 53116 70420 53172 71036
rect 53228 71026 53284 71036
rect 54124 71090 54180 72268
rect 54124 71038 54126 71090
rect 54178 71038 54180 71090
rect 54124 71026 54180 71038
rect 54236 70644 54292 73892
rect 54460 73892 54516 75292
rect 54796 75236 54852 75246
rect 54796 75122 54852 75180
rect 54796 75070 54798 75122
rect 54850 75070 54852 75122
rect 54796 75058 54852 75070
rect 54908 74900 54964 76524
rect 55020 76514 55076 76524
rect 55132 75684 55188 75694
rect 55132 75590 55188 75628
rect 55020 75460 55076 75470
rect 55020 75366 55076 75404
rect 55244 75458 55300 75470
rect 55244 75406 55246 75458
rect 55298 75406 55300 75458
rect 54796 74844 54964 74900
rect 55020 75236 55076 75246
rect 54460 73108 54516 73836
rect 54572 74340 54628 74350
rect 54572 73554 54628 74284
rect 54684 74116 54740 74126
rect 54684 74022 54740 74060
rect 54572 73502 54574 73554
rect 54626 73502 54628 73554
rect 54572 73490 54628 73502
rect 54460 73052 54628 73108
rect 54460 72772 54516 72782
rect 54348 72436 54404 72446
rect 54348 72342 54404 72380
rect 54460 71986 54516 72716
rect 54460 71934 54462 71986
rect 54514 71934 54516 71986
rect 54460 71202 54516 71934
rect 54460 71150 54462 71202
rect 54514 71150 54516 71202
rect 54460 71090 54516 71150
rect 54460 71038 54462 71090
rect 54514 71038 54516 71090
rect 54460 71026 54516 71038
rect 53060 70364 53172 70420
rect 54124 70588 54292 70644
rect 53004 70288 53060 70364
rect 54124 70308 54180 70588
rect 54572 70532 54628 73052
rect 54684 72548 54740 72558
rect 54684 72454 54740 72492
rect 54572 70466 54628 70476
rect 54684 71202 54740 71214
rect 54684 71150 54686 71202
rect 54738 71150 54740 71202
rect 54236 70420 54292 70430
rect 54236 70326 54292 70364
rect 54684 70418 54740 71150
rect 54684 70366 54686 70418
rect 54738 70366 54740 70418
rect 54684 70354 54740 70366
rect 54124 70242 54180 70252
rect 53452 70084 53508 70094
rect 53452 69990 53508 70028
rect 44716 69970 44772 69982
rect 44716 69918 44718 69970
rect 44770 69918 44772 69970
rect 44492 69524 44548 69534
rect 44380 69522 44548 69524
rect 44380 69470 44494 69522
rect 44546 69470 44548 69522
rect 44380 69468 44548 69470
rect 44716 69524 44772 69918
rect 44828 69524 44884 69534
rect 44716 69522 44884 69524
rect 44716 69470 44830 69522
rect 44882 69470 44884 69522
rect 44716 69468 44884 69470
rect 44492 69458 44548 69468
rect 44828 69458 44884 69468
rect 54684 69524 54740 69534
rect 54796 69524 54852 74844
rect 55020 74114 55076 75180
rect 55244 75236 55300 75406
rect 55244 75170 55300 75180
rect 55356 75124 55412 79200
rect 55356 75058 55412 75068
rect 55580 75682 55636 75694
rect 55580 75630 55582 75682
rect 55634 75630 55636 75682
rect 55580 75572 55636 75630
rect 55020 74062 55022 74114
rect 55074 74062 55076 74114
rect 55020 74050 55076 74062
rect 55244 74674 55300 74686
rect 55244 74622 55246 74674
rect 55298 74622 55300 74674
rect 54908 73892 54964 73902
rect 54908 73798 54964 73836
rect 54908 73444 54964 73454
rect 54908 73350 54964 73388
rect 54908 72772 54964 72782
rect 54908 72658 54964 72716
rect 54908 72606 54910 72658
rect 54962 72606 54964 72658
rect 54908 72594 54964 72606
rect 55244 71876 55300 74622
rect 55468 74676 55524 74686
rect 55356 73892 55412 73902
rect 55356 73556 55412 73836
rect 55356 73424 55412 73500
rect 55468 72436 55524 74620
rect 55580 72770 55636 75516
rect 56028 75348 56084 79200
rect 56588 77588 56644 77598
rect 56140 76354 56196 76366
rect 56140 76302 56142 76354
rect 56194 76302 56196 76354
rect 56140 75908 56196 76302
rect 56364 75908 56420 75918
rect 56196 75852 56308 75908
rect 56140 75842 56196 75852
rect 56140 75460 56196 75470
rect 56140 75366 56196 75404
rect 56028 75282 56084 75292
rect 55804 75236 55860 75246
rect 55692 74900 55748 74910
rect 55692 74786 55748 74844
rect 55692 74734 55694 74786
rect 55746 74734 55748 74786
rect 55692 74340 55748 74734
rect 55692 74274 55748 74284
rect 55692 74116 55748 74126
rect 55804 74116 55860 75180
rect 55692 74114 55972 74116
rect 55692 74062 55694 74114
rect 55746 74062 55972 74114
rect 55692 74060 55972 74062
rect 55692 74050 55748 74060
rect 55804 73890 55860 73902
rect 55804 73838 55806 73890
rect 55858 73838 55860 73890
rect 55580 72718 55582 72770
rect 55634 72718 55636 72770
rect 55580 72706 55636 72718
rect 55692 73220 55748 73230
rect 55692 72546 55748 73164
rect 55804 73108 55860 73838
rect 55916 73554 55972 74060
rect 56028 74004 56084 74042
rect 56028 73938 56084 73948
rect 55916 73502 55918 73554
rect 55970 73502 55972 73554
rect 55916 73444 55972 73502
rect 56028 73556 56084 73566
rect 56028 73462 56084 73500
rect 55916 73378 55972 73388
rect 56140 73332 56196 73342
rect 56028 73330 56196 73332
rect 56028 73278 56142 73330
rect 56194 73278 56196 73330
rect 56028 73276 56196 73278
rect 56028 73108 56084 73276
rect 56140 73266 56196 73276
rect 56252 73220 56308 75852
rect 56364 73332 56420 75852
rect 56476 75572 56532 75582
rect 56476 75478 56532 75516
rect 56588 75122 56644 77532
rect 56700 76580 56756 79200
rect 57372 76580 57428 79200
rect 56700 76514 56756 76524
rect 57148 76524 57428 76580
rect 57932 76580 57988 76590
rect 56924 76354 56980 76366
rect 56924 76302 56926 76354
rect 56978 76302 56980 76354
rect 56924 75908 56980 76302
rect 56924 75842 56980 75852
rect 57036 75458 57092 75470
rect 57036 75406 57038 75458
rect 57090 75406 57092 75458
rect 57036 75236 57092 75406
rect 57036 75170 57092 75180
rect 56588 75070 56590 75122
rect 56642 75070 56644 75122
rect 56588 75058 56644 75070
rect 56924 74674 56980 74686
rect 56924 74622 56926 74674
rect 56978 74622 56980 74674
rect 56588 74228 56644 74238
rect 56588 73556 56644 74172
rect 56924 74116 56980 74622
rect 56924 74050 56980 74060
rect 57036 74676 57092 74686
rect 56812 74002 56868 74014
rect 56812 73950 56814 74002
rect 56866 73950 56868 74002
rect 56588 73500 56756 73556
rect 56588 73332 56644 73342
rect 56364 73330 56644 73332
rect 56364 73278 56590 73330
rect 56642 73278 56644 73330
rect 56364 73276 56644 73278
rect 56252 73154 56308 73164
rect 55804 73052 56084 73108
rect 55692 72494 55694 72546
rect 55746 72494 55748 72546
rect 55692 72482 55748 72494
rect 55580 72436 55636 72446
rect 55468 72434 55636 72436
rect 55468 72382 55582 72434
rect 55634 72382 55636 72434
rect 55468 72380 55636 72382
rect 55244 71762 55300 71820
rect 55244 71710 55246 71762
rect 55298 71710 55300 71762
rect 54908 71202 54964 71214
rect 54908 71150 54910 71202
rect 54962 71150 54964 71202
rect 54908 71090 54964 71150
rect 54908 71038 54910 71090
rect 54962 71038 54964 71090
rect 54908 71026 54964 71038
rect 55244 70756 55300 71710
rect 55468 71874 55524 71886
rect 55468 71822 55470 71874
rect 55522 71822 55524 71874
rect 55468 70980 55524 71822
rect 55468 70914 55524 70924
rect 55244 70690 55300 70700
rect 55468 70756 55524 70766
rect 55468 70662 55524 70700
rect 55356 70532 55412 70542
rect 55356 70418 55412 70476
rect 55356 70366 55358 70418
rect 55410 70366 55412 70418
rect 55356 70354 55412 70366
rect 55580 70420 55636 72380
rect 55916 70980 55972 70990
rect 56028 70980 56084 73052
rect 56588 73108 56644 73276
rect 56588 73042 56644 73052
rect 56476 72658 56532 72670
rect 56476 72606 56478 72658
rect 56530 72606 56532 72658
rect 56140 71204 56196 71214
rect 56140 71110 56196 71148
rect 56476 71202 56532 72606
rect 56700 72324 56756 73500
rect 56812 73220 56868 73950
rect 57036 74002 57092 74620
rect 57036 73950 57038 74002
rect 57090 73950 57092 74002
rect 57036 73938 57092 73950
rect 56924 73890 56980 73902
rect 56924 73838 56926 73890
rect 56978 73838 56980 73890
rect 56924 73332 56980 73838
rect 57148 73892 57204 76524
rect 57932 76486 57988 76524
rect 57372 75570 57428 75582
rect 57372 75518 57374 75570
rect 57426 75518 57428 75570
rect 57372 75236 57428 75518
rect 57932 75460 57988 75470
rect 57372 75170 57428 75180
rect 57708 75458 57988 75460
rect 57708 75406 57934 75458
rect 57986 75406 57988 75458
rect 57708 75404 57988 75406
rect 57484 75012 57540 75022
rect 57148 73826 57204 73836
rect 57260 75010 57540 75012
rect 57260 74958 57486 75010
rect 57538 74958 57540 75010
rect 57260 74956 57540 74958
rect 57260 73442 57316 74956
rect 57484 74946 57540 74956
rect 57708 74898 57764 75404
rect 57932 75394 57988 75404
rect 58044 75460 58100 79200
rect 58716 76804 58772 79200
rect 59388 76804 59444 79200
rect 60060 76916 60116 79200
rect 60620 77364 60676 77374
rect 60060 76860 60228 76916
rect 58716 76748 59220 76804
rect 59388 76748 60116 76804
rect 58604 76580 58660 76590
rect 58380 76132 58436 76142
rect 58044 75394 58100 75404
rect 58268 75458 58324 75470
rect 58268 75406 58270 75458
rect 58322 75406 58324 75458
rect 57708 74846 57710 74898
rect 57762 74846 57764 74898
rect 57596 74116 57652 74126
rect 57596 74022 57652 74060
rect 57708 73948 57764 74846
rect 58044 75236 58100 75246
rect 57260 73390 57262 73442
rect 57314 73390 57316 73442
rect 57260 73378 57316 73390
rect 57484 73892 57764 73948
rect 57932 74004 57988 74042
rect 57932 73938 57988 73948
rect 57484 73780 57540 73892
rect 56924 73266 56980 73276
rect 56812 73154 56868 73164
rect 57148 72770 57204 72782
rect 57148 72718 57150 72770
rect 57202 72718 57204 72770
rect 57148 72660 57204 72718
rect 57148 72594 57204 72604
rect 57484 72660 57540 73724
rect 57820 73890 57876 73902
rect 57820 73838 57822 73890
rect 57874 73838 57876 73890
rect 57820 73556 57876 73838
rect 57820 73490 57876 73500
rect 58044 73444 58100 75180
rect 58268 75012 58324 75406
rect 58268 74946 58324 74956
rect 58268 74788 58324 74798
rect 58380 74788 58436 76076
rect 58268 74786 58436 74788
rect 58268 74734 58270 74786
rect 58322 74734 58436 74786
rect 58268 74732 58436 74734
rect 58268 74564 58324 74732
rect 58268 74498 58324 74508
rect 58604 73780 58660 76524
rect 58940 76578 58996 76590
rect 58940 76526 58942 76578
rect 58994 76526 58996 76578
rect 58940 75796 58996 76526
rect 59164 76468 59220 76748
rect 59836 76578 59892 76590
rect 59836 76526 59838 76578
rect 59890 76526 59892 76578
rect 59836 76468 59892 76526
rect 59164 76466 59556 76468
rect 59164 76414 59166 76466
rect 59218 76414 59556 76466
rect 59164 76412 59556 76414
rect 59164 76402 59220 76412
rect 58940 75730 58996 75740
rect 59164 75908 59220 75918
rect 59164 75570 59220 75852
rect 59164 75518 59166 75570
rect 59218 75518 59220 75570
rect 58828 75460 58884 75470
rect 58828 75458 58996 75460
rect 58828 75406 58830 75458
rect 58882 75406 58996 75458
rect 58828 75404 58996 75406
rect 58828 75394 58884 75404
rect 58940 75124 58996 75404
rect 59164 75124 59220 75518
rect 59500 75236 59556 76412
rect 59836 76402 59892 76412
rect 59612 76020 59668 76030
rect 59612 75682 59668 75964
rect 59612 75630 59614 75682
rect 59666 75630 59668 75682
rect 59612 75618 59668 75630
rect 59948 75572 60004 75582
rect 59836 75458 59892 75470
rect 59836 75406 59838 75458
rect 59890 75406 59892 75458
rect 59836 75236 59892 75406
rect 59500 75180 59668 75236
rect 59276 75124 59332 75134
rect 59164 75122 59332 75124
rect 59164 75070 59278 75122
rect 59330 75070 59332 75122
rect 59164 75068 59332 75070
rect 58940 75058 58996 75068
rect 58828 75012 58884 75022
rect 58828 74898 58884 74956
rect 59164 74900 59220 74910
rect 58828 74846 58830 74898
rect 58882 74846 58884 74898
rect 58828 74788 58884 74846
rect 58716 74116 58772 74126
rect 58828 74116 58884 74732
rect 58716 74114 58884 74116
rect 58716 74062 58718 74114
rect 58770 74062 58884 74114
rect 58716 74060 58884 74062
rect 58940 74844 59164 74900
rect 58940 74114 58996 74844
rect 59164 74806 59220 74844
rect 58940 74062 58942 74114
rect 58994 74062 58996 74114
rect 58716 74050 58772 74060
rect 58940 74050 58996 74062
rect 59164 74228 59220 74238
rect 58828 73892 58884 73902
rect 58828 73890 58996 73892
rect 58828 73838 58830 73890
rect 58882 73838 58996 73890
rect 58828 73836 58996 73838
rect 58828 73826 58884 73836
rect 58604 73714 58660 73724
rect 58044 73388 58212 73444
rect 57708 73332 57764 73342
rect 57764 73276 57988 73332
rect 57708 73238 57764 73276
rect 57484 72594 57540 72604
rect 56476 71150 56478 71202
rect 56530 71150 56532 71202
rect 56476 71138 56532 71150
rect 56588 72268 56756 72324
rect 57036 72546 57092 72558
rect 57036 72494 57038 72546
rect 57090 72494 57092 72546
rect 57036 72436 57092 72494
rect 55972 70924 56084 70980
rect 55916 70886 55972 70924
rect 55580 70084 55636 70364
rect 56028 70420 56084 70430
rect 56028 70326 56084 70364
rect 56476 70420 56532 70430
rect 56476 70326 56532 70364
rect 56588 70308 56644 72268
rect 56700 72100 56756 72110
rect 56700 71876 56756 72044
rect 56700 71744 56756 71820
rect 56924 71764 56980 71774
rect 57036 71764 57092 72380
rect 56924 71762 57092 71764
rect 56924 71710 56926 71762
rect 56978 71710 57092 71762
rect 56924 71708 57092 71710
rect 57260 72546 57316 72558
rect 57260 72494 57262 72546
rect 57314 72494 57316 72546
rect 56924 71698 56980 71708
rect 57260 71090 57316 72494
rect 57932 72546 57988 73276
rect 57932 72494 57934 72546
rect 57986 72494 57988 72546
rect 57932 72482 57988 72494
rect 58044 73218 58100 73230
rect 58044 73166 58046 73218
rect 58098 73166 58100 73218
rect 58044 72658 58100 73166
rect 58044 72606 58046 72658
rect 58098 72606 58100 72658
rect 58044 71986 58100 72606
rect 58044 71934 58046 71986
rect 58098 71934 58100 71986
rect 58044 71922 58100 71934
rect 57260 71038 57262 71090
rect 57314 71038 57316 71090
rect 57372 71876 57428 71886
rect 57372 71204 57428 71820
rect 57932 71876 57988 71886
rect 57932 71782 57988 71820
rect 57372 71072 57428 71148
rect 57932 71092 57988 71102
rect 58156 71092 58212 73388
rect 58828 73218 58884 73230
rect 58828 73166 58830 73218
rect 58882 73166 58884 73218
rect 58828 72548 58884 73166
rect 58828 72482 58884 72492
rect 58716 72100 58772 72110
rect 58716 71986 58772 72044
rect 58716 71934 58718 71986
rect 58770 71934 58772 71986
rect 58716 71922 58772 71934
rect 58940 71876 58996 73836
rect 59164 73332 59220 74172
rect 59276 74114 59332 75068
rect 59500 74898 59556 74910
rect 59500 74846 59502 74898
rect 59554 74846 59556 74898
rect 59276 74062 59278 74114
rect 59330 74062 59332 74114
rect 59276 74050 59332 74062
rect 59388 74786 59444 74798
rect 59388 74734 59390 74786
rect 59442 74734 59444 74786
rect 59276 73332 59332 73370
rect 59164 73276 59276 73332
rect 59276 73266 59332 73276
rect 59388 73220 59444 74734
rect 59500 74340 59556 74846
rect 59500 74274 59556 74284
rect 59612 73444 59668 75180
rect 59836 75170 59892 75180
rect 59724 75012 59780 75022
rect 59724 74564 59780 74956
rect 59948 75012 60004 75516
rect 59948 74946 60004 74956
rect 59724 74498 59780 74508
rect 60060 73948 60116 76748
rect 60172 75236 60228 76860
rect 60508 76692 60564 76702
rect 60508 76598 60564 76636
rect 60508 75572 60564 75582
rect 60620 75572 60676 77308
rect 60732 77026 60788 79200
rect 60732 76974 60734 77026
rect 60786 76974 60788 77026
rect 60732 76962 60788 76974
rect 60508 75570 60676 75572
rect 60508 75518 60510 75570
rect 60562 75518 60676 75570
rect 60508 75516 60676 75518
rect 61404 75572 61460 79200
rect 61964 77026 62020 77038
rect 61964 76974 61966 77026
rect 62018 76974 62020 77026
rect 61964 76690 62020 76974
rect 61964 76638 61966 76690
rect 62018 76638 62020 76690
rect 61628 76578 61684 76590
rect 61628 76526 61630 76578
rect 61682 76526 61684 76578
rect 61628 75684 61684 76526
rect 61628 75618 61684 75628
rect 60508 75506 60564 75516
rect 61404 75506 61460 75516
rect 61740 75458 61796 75470
rect 61740 75406 61742 75458
rect 61794 75406 61796 75458
rect 61740 75348 61796 75406
rect 61740 75282 61796 75292
rect 60172 75170 60228 75180
rect 61628 75124 61684 75134
rect 60172 75012 60228 75022
rect 60172 74918 60228 74956
rect 61628 75012 61684 75068
rect 61852 75012 61908 75022
rect 61628 75010 61852 75012
rect 61628 74958 61630 75010
rect 61682 74958 61852 75010
rect 61628 74956 61852 74958
rect 61628 74946 61684 74956
rect 61516 74900 61572 74910
rect 61516 74806 61572 74844
rect 60284 74788 60340 74798
rect 60284 74694 60340 74732
rect 60956 74786 61012 74798
rect 60956 74734 60958 74786
rect 61010 74734 61012 74786
rect 60844 74676 60900 74686
rect 60844 74582 60900 74620
rect 60956 74564 61012 74734
rect 60956 74498 61012 74508
rect 61404 74788 61460 74798
rect 60620 74340 60676 74350
rect 59836 73890 59892 73902
rect 60060 73892 60228 73948
rect 59836 73838 59838 73890
rect 59890 73838 59892 73890
rect 59836 73668 59892 73838
rect 60172 73780 60228 73892
rect 60508 73892 60564 73902
rect 60508 73798 60564 73836
rect 60172 73724 60452 73780
rect 59836 73602 59892 73612
rect 60396 73554 60452 73724
rect 60396 73502 60398 73554
rect 60450 73502 60452 73554
rect 60396 73490 60452 73502
rect 59612 73388 59780 73444
rect 59612 73220 59668 73230
rect 59388 73218 59668 73220
rect 59388 73166 59614 73218
rect 59666 73166 59668 73218
rect 59388 73164 59668 73166
rect 59612 73154 59668 73164
rect 59276 73108 59332 73118
rect 59276 72658 59332 73052
rect 59724 72996 59780 73388
rect 59276 72606 59278 72658
rect 59330 72606 59332 72658
rect 59276 72594 59332 72606
rect 59612 72940 59780 72996
rect 60172 73332 60228 73342
rect 59164 72436 59220 72446
rect 59164 72342 59220 72380
rect 59276 71988 59332 71998
rect 59276 71894 59332 71932
rect 59612 71986 59668 72940
rect 59724 72660 59780 72670
rect 59724 72566 59780 72604
rect 60172 72658 60228 73276
rect 60620 72660 60676 74284
rect 61404 74116 61460 74732
rect 61628 74340 61684 74350
rect 61628 74226 61684 74284
rect 61628 74174 61630 74226
rect 61682 74174 61684 74226
rect 61628 74162 61684 74174
rect 60956 73780 61012 73790
rect 60956 73554 61012 73724
rect 60956 73502 60958 73554
rect 61010 73502 61012 73554
rect 60956 73490 61012 73502
rect 61404 73554 61460 74060
rect 61404 73502 61406 73554
rect 61458 73502 61460 73554
rect 60172 72606 60174 72658
rect 60226 72606 60228 72658
rect 60172 72594 60228 72606
rect 60396 72658 60676 72660
rect 60396 72606 60622 72658
rect 60674 72606 60676 72658
rect 60396 72604 60676 72606
rect 60396 72100 60452 72604
rect 60620 72594 60676 72604
rect 60396 72034 60452 72044
rect 59612 71934 59614 71986
rect 59666 71934 59668 71986
rect 59612 71922 59668 71934
rect 61404 71988 61460 73502
rect 61852 73554 61908 74956
rect 61964 74228 62020 76638
rect 62076 75124 62132 79200
rect 62748 76580 62804 79200
rect 63420 77364 63476 79200
rect 63420 77308 63812 77364
rect 62748 76514 62804 76524
rect 63532 76580 63588 76590
rect 62412 76468 62468 76478
rect 62412 76374 62468 76412
rect 62860 76244 62916 76254
rect 62860 76150 62916 76188
rect 62524 76132 62580 76142
rect 62412 75460 62468 75470
rect 62412 75366 62468 75404
rect 62076 75058 62132 75068
rect 62188 75236 62244 75246
rect 62188 75122 62244 75180
rect 62188 75070 62190 75122
rect 62242 75070 62244 75122
rect 62188 75058 62244 75070
rect 62524 74228 62580 76076
rect 63084 75572 63140 75582
rect 63084 75478 63140 75516
rect 62860 75124 62916 75134
rect 62860 75030 62916 75068
rect 63420 74788 63476 74798
rect 63420 74694 63476 74732
rect 61964 74162 62020 74172
rect 62076 74226 62580 74228
rect 62076 74174 62526 74226
rect 62578 74174 62580 74226
rect 62076 74172 62580 74174
rect 62076 74116 62132 74172
rect 62524 74162 62580 74172
rect 62972 74228 63028 74238
rect 62972 74134 63028 74172
rect 63532 74226 63588 76524
rect 63756 75570 63812 77308
rect 63756 75518 63758 75570
rect 63810 75518 63812 75570
rect 63756 75506 63812 75518
rect 63868 75572 63924 75582
rect 64092 75572 64148 79200
rect 64764 77140 64820 79200
rect 64764 77084 65268 77140
rect 64988 76580 65044 76590
rect 64988 76486 65044 76524
rect 65212 76580 65268 77084
rect 65212 75794 65268 76524
rect 65212 75742 65214 75794
rect 65266 75742 65268 75794
rect 65212 75730 65268 75742
rect 64428 75572 64484 75582
rect 64092 75570 64484 75572
rect 64092 75518 64430 75570
rect 64482 75518 64484 75570
rect 64092 75516 64484 75518
rect 65436 75572 65492 79200
rect 66108 77364 66164 79200
rect 66108 77308 66388 77364
rect 65884 76244 65940 76254
rect 65772 76242 65940 76244
rect 65772 76190 65886 76242
rect 65938 76190 65940 76242
rect 65772 76188 65940 76190
rect 65660 75572 65716 75582
rect 65436 75570 65716 75572
rect 65436 75518 65662 75570
rect 65714 75518 65716 75570
rect 65436 75516 65716 75518
rect 63868 75122 63924 75516
rect 64428 75506 64484 75516
rect 65660 75506 65716 75516
rect 63868 75070 63870 75122
rect 63922 75070 63924 75122
rect 63868 75012 63924 75070
rect 63868 74946 63924 74956
rect 65772 74340 65828 76188
rect 65884 76178 65940 76188
rect 65916 76076 66180 76086
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 65916 76010 66180 76020
rect 66332 75570 66388 77308
rect 66332 75518 66334 75570
rect 66386 75518 66388 75570
rect 66332 75506 66388 75518
rect 66780 75572 66836 79200
rect 67452 77140 67508 79200
rect 67452 77084 67732 77140
rect 66780 75122 66836 75516
rect 66780 75070 66782 75122
rect 66834 75070 66836 75122
rect 66780 75058 66836 75070
rect 66892 75458 66948 75470
rect 66892 75406 66894 75458
rect 66946 75406 66948 75458
rect 65916 74508 66180 74518
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 65916 74442 66180 74452
rect 65772 74274 65828 74284
rect 63532 74174 63534 74226
rect 63586 74174 63588 74226
rect 63532 74162 63588 74174
rect 62076 74022 62132 74060
rect 61852 73502 61854 73554
rect 61906 73502 61908 73554
rect 61852 73490 61908 73502
rect 66892 73332 66948 75406
rect 67676 75122 67732 77084
rect 68124 76692 68180 79200
rect 68796 76804 68852 79200
rect 68796 76738 68852 76748
rect 69356 76804 69412 76814
rect 68124 76626 68180 76636
rect 69356 76690 69412 76748
rect 69356 76638 69358 76690
rect 69410 76638 69412 76690
rect 69356 76626 69412 76638
rect 68012 76580 68068 76590
rect 68012 76486 68068 76524
rect 69020 76578 69076 76590
rect 69020 76526 69022 76578
rect 69074 76526 69076 76578
rect 69020 76356 69076 76526
rect 69020 76290 69076 76300
rect 69020 75572 69076 75582
rect 69020 75478 69076 75516
rect 69468 75460 69524 79200
rect 69916 76692 69972 76702
rect 69916 76598 69972 76636
rect 70140 75572 70196 79200
rect 70476 76804 70532 76814
rect 70476 76690 70532 76748
rect 70476 76638 70478 76690
rect 70530 76638 70532 76690
rect 70476 76626 70532 76638
rect 70812 76580 70868 79200
rect 70924 77476 70980 77486
rect 70924 76690 70980 77420
rect 70924 76638 70926 76690
rect 70978 76638 70980 76690
rect 70924 76626 70980 76638
rect 70140 75506 70196 75516
rect 70700 75572 70756 75582
rect 70700 75478 70756 75516
rect 69468 75394 69524 75404
rect 70028 75460 70084 75470
rect 70028 75366 70084 75404
rect 67676 75070 67678 75122
rect 67730 75070 67732 75122
rect 67676 75058 67732 75070
rect 70812 75122 70868 76524
rect 71484 75572 71540 79200
rect 71708 75572 71764 75582
rect 71484 75570 71764 75572
rect 71484 75518 71710 75570
rect 71762 75518 71764 75570
rect 71484 75516 71764 75518
rect 72156 75572 72212 79200
rect 72380 75572 72436 75582
rect 72156 75570 72436 75572
rect 72156 75518 72382 75570
rect 72434 75518 72436 75570
rect 72156 75516 72436 75518
rect 71708 75506 71764 75516
rect 72380 75506 72436 75516
rect 70812 75070 70814 75122
rect 70866 75070 70868 75122
rect 70812 75058 70868 75070
rect 72828 75460 72884 79200
rect 73052 76580 73108 76590
rect 73052 76486 73108 76524
rect 73388 75570 73444 75582
rect 73388 75518 73390 75570
rect 73442 75518 73444 75570
rect 72828 75122 72884 75404
rect 72828 75070 72830 75122
rect 72882 75070 72884 75122
rect 72828 75058 72884 75070
rect 73052 75458 73108 75470
rect 73052 75406 73054 75458
rect 73106 75406 73108 75458
rect 66892 73266 66948 73276
rect 65916 72940 66180 72950
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 65916 72874 66180 72884
rect 61404 71922 61460 71932
rect 58940 71810 58996 71820
rect 65916 71372 66180 71382
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 65916 71306 66180 71316
rect 57932 71090 58212 71092
rect 57260 71026 57316 71038
rect 57932 71038 57934 71090
rect 57986 71038 58212 71090
rect 57932 71036 58212 71038
rect 73052 71092 73108 75406
rect 73388 75460 73444 75518
rect 73500 75572 73556 79200
rect 73500 75506 73556 75516
rect 73948 75572 74004 75582
rect 73948 75478 74004 75516
rect 73388 75394 73444 75404
rect 74172 75124 74228 79200
rect 74508 76244 74564 76254
rect 74508 76150 74564 76188
rect 74844 75684 74900 79200
rect 75068 75794 75124 75806
rect 75068 75742 75070 75794
rect 75122 75742 75124 75794
rect 75068 75684 75124 75742
rect 74844 75628 75012 75684
rect 74956 75572 75012 75628
rect 75068 75618 75124 75628
rect 75516 75572 75572 79200
rect 76188 77140 76244 79200
rect 76188 77084 76468 77140
rect 75516 75516 75796 75572
rect 74956 75506 75012 75516
rect 74396 75124 74452 75134
rect 74172 75122 74452 75124
rect 74172 75070 74398 75122
rect 74450 75070 74452 75122
rect 74172 75068 74452 75070
rect 74396 75058 74452 75068
rect 75740 75122 75796 75516
rect 75740 75070 75742 75122
rect 75794 75070 75796 75122
rect 75740 75058 75796 75070
rect 76412 75122 76468 77084
rect 76860 76580 76916 79200
rect 77532 77364 77588 79200
rect 77532 77308 78036 77364
rect 77644 76580 77700 76590
rect 76860 76578 77700 76580
rect 76860 76526 77646 76578
rect 77698 76526 77700 76578
rect 76860 76524 77700 76526
rect 76972 75572 77028 75582
rect 76972 75478 77028 75516
rect 77420 75572 77476 75582
rect 76412 75070 76414 75122
rect 76466 75070 76468 75122
rect 76412 75058 76468 75070
rect 77420 75122 77476 75516
rect 77420 75070 77422 75122
rect 77474 75070 77476 75122
rect 77420 75058 77476 75070
rect 77644 74228 77700 76524
rect 77980 75570 78036 77308
rect 77980 75518 77982 75570
rect 78034 75518 78036 75570
rect 77980 75506 78036 75518
rect 78092 75124 78148 75134
rect 78204 75124 78260 79200
rect 78092 75122 78260 75124
rect 78092 75070 78094 75122
rect 78146 75070 78260 75122
rect 78092 75068 78260 75070
rect 78092 75058 78148 75068
rect 77644 74162 77700 74172
rect 78092 74228 78148 74238
rect 78092 74134 78148 74172
rect 57932 71026 57988 71036
rect 73052 71026 73108 71036
rect 57036 70980 57092 70990
rect 57036 70886 57092 70924
rect 56588 70242 56644 70252
rect 56924 70308 56980 70318
rect 56924 70214 56980 70252
rect 55580 70018 55636 70028
rect 65916 69804 66180 69814
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 65916 69738 66180 69748
rect 54684 69522 54852 69524
rect 54684 69470 54686 69522
rect 54738 69470 54852 69522
rect 54684 69468 54852 69470
rect 54684 69458 54740 69468
rect 19836 69020 20100 69030
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 19836 68954 20100 68964
rect 50556 69020 50820 69030
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50556 68954 50820 68964
rect 4476 68236 4740 68246
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4476 68170 4740 68180
rect 35196 68236 35460 68246
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35196 68170 35460 68180
rect 65916 68236 66180 68246
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 65916 68170 66180 68180
rect 19836 67452 20100 67462
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 19836 67386 20100 67396
rect 50556 67452 50820 67462
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50556 67386 50820 67396
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 35196 66668 35460 66678
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35196 66602 35460 66612
rect 65916 66668 66180 66678
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 65916 66602 66180 66612
rect 19836 65884 20100 65894
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 19836 65818 20100 65828
rect 50556 65884 50820 65894
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50556 65818 50820 65828
rect 4476 65100 4740 65110
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 35196 65100 35460 65110
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35196 65034 35460 65044
rect 65916 65100 66180 65110
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 65916 65034 66180 65044
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 50556 64316 50820 64326
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50556 64250 50820 64260
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35196 63466 35460 63476
rect 65916 63532 66180 63542
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 65916 63466 66180 63476
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 50556 62748 50820 62758
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50556 62682 50820 62692
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 65916 61964 66180 61974
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 65916 61898 66180 61908
rect 19836 61180 20100 61190
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 50556 61180 50820 61190
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50556 61114 50820 61124
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 65916 60396 66180 60406
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 65916 60330 66180 60340
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 50556 59612 50820 59622
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50556 59546 50820 59556
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 65916 58828 66180 58838
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 65916 58762 66180 58772
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 50556 58044 50820 58054
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50556 57978 50820 57988
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 65916 57260 66180 57270
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 65916 57194 66180 57204
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 65916 55692 66180 55702
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 65916 55626 66180 55636
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 65916 54124 66180 54134
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 65916 54058 66180 54068
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 65916 52556 66180 52566
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 65916 52490 66180 52500
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 65916 50988 66180 50998
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 65916 50922 66180 50932
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 65916 49420 66180 49430
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 65916 49354 66180 49364
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 65916 47852 66180 47862
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 65916 47786 66180 47796
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 65916 46284 66180 46294
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 65916 46218 66180 46228
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 65916 44716 66180 44726
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 65916 44650 66180 44660
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 65916 43148 66180 43158
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 65916 43082 66180 43092
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 65916 41580 66180 41590
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 65916 41514 66180 41524
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 65916 40012 66180 40022
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 65916 39946 66180 39956
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 65916 38444 66180 38454
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 65916 38378 66180 38388
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 65916 36876 66180 36886
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 65916 36810 66180 36820
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 65916 35308 66180 35318
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 65916 35242 66180 35252
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 65916 33740 66180 33750
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 65916 33674 66180 33684
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 65916 32172 66180 32182
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 65916 32106 66180 32116
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 65916 30604 66180 30614
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 65916 30538 66180 30548
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 65916 29036 66180 29046
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 65916 28970 66180 28980
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 65916 27468 66180 27478
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 65916 27402 66180 27412
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 65916 25900 66180 25910
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 65916 25834 66180 25844
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 65916 24332 66180 24342
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 65916 24266 66180 24276
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 65916 22764 66180 22774
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 65916 22698 66180 22708
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 65916 21196 66180 21206
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 65916 21130 66180 21140
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 65916 19628 66180 19638
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 65916 19562 66180 19572
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 65916 18060 66180 18070
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 65916 17994 66180 18004
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 65916 16492 66180 16502
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 65916 16426 66180 16436
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 65916 14924 66180 14934
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 65916 14858 66180 14868
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 65916 13356 66180 13366
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 65916 13290 66180 13300
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 65916 11788 66180 11798
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 65916 11722 66180 11732
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 65916 10220 66180 10230
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 65916 10154 66180 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 65916 8652 66180 8662
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 65916 8586 66180 8596
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 65916 7084 66180 7094
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 65916 7018 66180 7028
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 65916 5516 66180 5526
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 65916 5450 66180 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 73276 4452 73332 4462
rect 73948 4452 74004 4462
rect 73164 4450 73332 4452
rect 73164 4398 73278 4450
rect 73330 4398 73332 4450
rect 73164 4396 73332 4398
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 65916 3948 66180 3958
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 65916 3882 66180 3892
rect 6972 3332 7028 3342
rect 8316 3332 8372 3342
rect 9212 3332 9268 3342
rect 10108 3332 10164 3342
rect 6748 3330 7028 3332
rect 6748 3278 6974 3330
rect 7026 3278 7028 3330
rect 6748 3276 7028 3278
rect 6748 800 6804 3276
rect 6972 3266 7028 3276
rect 8092 3330 8372 3332
rect 8092 3278 8318 3330
rect 8370 3278 8372 3330
rect 8092 3276 8372 3278
rect 8092 800 8148 3276
rect 8316 3266 8372 3276
rect 8988 3330 9268 3332
rect 8988 3278 9214 3330
rect 9266 3278 9268 3330
rect 8988 3276 9268 3278
rect 8988 800 9044 3276
rect 9212 3266 9268 3276
rect 9884 3330 10164 3332
rect 9884 3278 10110 3330
rect 10162 3278 10164 3330
rect 9884 3276 10164 3278
rect 9884 800 9940 3276
rect 10108 3266 10164 3276
rect 10780 3330 10836 3342
rect 10780 3278 10782 3330
rect 10834 3278 10836 3330
rect 10780 800 10836 3278
rect 11564 3332 11620 3342
rect 12236 3332 12292 3342
rect 12908 3332 12964 3342
rect 13580 3332 13636 3342
rect 14252 3332 14308 3342
rect 14924 3332 14980 3342
rect 15596 3332 15652 3342
rect 16268 3332 16324 3342
rect 16940 3332 16996 3342
rect 17612 3332 17668 3342
rect 18284 3332 18340 3342
rect 18956 3332 19012 3342
rect 11564 3330 11732 3332
rect 11564 3278 11566 3330
rect 11618 3278 11732 3330
rect 11564 3276 11732 3278
rect 11564 3266 11620 3276
rect 11676 800 11732 3276
rect 12236 3330 12404 3332
rect 12236 3278 12238 3330
rect 12290 3278 12404 3330
rect 12236 3276 12404 3278
rect 12236 3266 12292 3276
rect 12348 800 12404 3276
rect 12908 3330 13076 3332
rect 12908 3278 12910 3330
rect 12962 3278 13076 3330
rect 12908 3276 13076 3278
rect 12908 3266 12964 3276
rect 13020 800 13076 3276
rect 13580 3330 13748 3332
rect 13580 3278 13582 3330
rect 13634 3278 13748 3330
rect 13580 3276 13748 3278
rect 13580 3266 13636 3276
rect 13692 800 13748 3276
rect 14252 3330 14420 3332
rect 14252 3278 14254 3330
rect 14306 3278 14420 3330
rect 14252 3276 14420 3278
rect 14252 3266 14308 3276
rect 14364 800 14420 3276
rect 14924 3330 15092 3332
rect 14924 3278 14926 3330
rect 14978 3278 15092 3330
rect 14924 3276 15092 3278
rect 14924 3266 14980 3276
rect 15036 800 15092 3276
rect 15596 3330 15764 3332
rect 15596 3278 15598 3330
rect 15650 3278 15764 3330
rect 15596 3276 15764 3278
rect 15596 3266 15652 3276
rect 15708 800 15764 3276
rect 16268 3330 16436 3332
rect 16268 3278 16270 3330
rect 16322 3278 16436 3330
rect 16268 3276 16436 3278
rect 16268 3266 16324 3276
rect 16380 800 16436 3276
rect 16940 3330 17108 3332
rect 16940 3278 16942 3330
rect 16994 3278 17108 3330
rect 16940 3276 17108 3278
rect 16940 3266 16996 3276
rect 17052 800 17108 3276
rect 17612 3330 17780 3332
rect 17612 3278 17614 3330
rect 17666 3278 17780 3330
rect 17612 3276 17780 3278
rect 17612 3266 17668 3276
rect 17724 800 17780 3276
rect 18284 3330 18452 3332
rect 18284 3278 18286 3330
rect 18338 3278 18452 3330
rect 18284 3276 18452 3278
rect 18284 3266 18340 3276
rect 18396 800 18452 3276
rect 18956 3330 19124 3332
rect 18956 3278 18958 3330
rect 19010 3278 19124 3330
rect 18956 3276 19124 3278
rect 18956 3266 19012 3276
rect 19068 800 19124 3276
rect 19628 3330 19684 3342
rect 19628 3278 19630 3330
rect 19682 3278 19684 3330
rect 19628 1652 19684 3278
rect 20300 3332 20356 3342
rect 20972 3332 21028 3342
rect 20300 3330 20468 3332
rect 20300 3278 20302 3330
rect 20354 3278 20468 3330
rect 20300 3276 20468 3278
rect 20300 3266 20356 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 19628 1596 19796 1652
rect 19740 800 19796 1596
rect 20412 800 20468 3276
rect 20972 3330 21140 3332
rect 20972 3278 20974 3330
rect 21026 3278 21140 3330
rect 20972 3276 21140 3278
rect 20972 3266 21028 3276
rect 21084 800 21140 3276
rect 21756 3330 21812 3342
rect 21756 3278 21758 3330
rect 21810 3278 21812 3330
rect 21756 800 21812 3278
rect 22428 3330 22484 3342
rect 22428 3278 22430 3330
rect 22482 3278 22484 3330
rect 22428 800 22484 3278
rect 23100 3330 23156 3342
rect 23100 3278 23102 3330
rect 23154 3278 23156 3330
rect 23100 800 23156 3278
rect 23772 3330 23828 3342
rect 23772 3278 23774 3330
rect 23826 3278 23828 3330
rect 23772 800 23828 3278
rect 24444 3330 24500 3342
rect 24444 3278 24446 3330
rect 24498 3278 24500 3330
rect 24444 800 24500 3278
rect 25116 3330 25172 3342
rect 25116 3278 25118 3330
rect 25170 3278 25172 3330
rect 25116 800 25172 3278
rect 25788 3330 25844 3342
rect 25788 3278 25790 3330
rect 25842 3278 25844 3330
rect 25788 800 25844 3278
rect 26460 3330 26516 3342
rect 26460 3278 26462 3330
rect 26514 3278 26516 3330
rect 26460 800 26516 3278
rect 27132 3330 27188 3342
rect 27132 3278 27134 3330
rect 27186 3278 27188 3330
rect 27132 800 27188 3278
rect 27804 3330 27860 3342
rect 27804 3278 27806 3330
rect 27858 3278 27860 3330
rect 27804 800 27860 3278
rect 28476 3330 28532 3342
rect 28476 3278 28478 3330
rect 28530 3278 28532 3330
rect 28476 800 28532 3278
rect 29148 3330 29204 3342
rect 29148 3278 29150 3330
rect 29202 3278 29204 3330
rect 29148 800 29204 3278
rect 29820 3330 29876 3342
rect 30492 3332 30548 3342
rect 31164 3332 31220 3342
rect 31836 3332 31892 3342
rect 32508 3332 32564 3342
rect 33180 3332 33236 3342
rect 33852 3332 33908 3342
rect 34524 3332 34580 3342
rect 35196 3332 35252 3342
rect 35868 3332 35924 3342
rect 36540 3332 36596 3342
rect 37212 3332 37268 3342
rect 37884 3332 37940 3342
rect 38556 3332 38612 3342
rect 39228 3332 39284 3342
rect 39900 3332 39956 3342
rect 40572 3332 40628 3342
rect 29820 3278 29822 3330
rect 29874 3278 29876 3330
rect 29820 800 29876 3278
rect 30268 3330 30548 3332
rect 30268 3278 30494 3330
rect 30546 3278 30548 3330
rect 30268 3276 30548 3278
rect 30268 800 30324 3276
rect 30492 3266 30548 3276
rect 30940 3330 31220 3332
rect 30940 3278 31166 3330
rect 31218 3278 31220 3330
rect 30940 3276 31220 3278
rect 30940 800 30996 3276
rect 31164 3266 31220 3276
rect 31612 3330 31892 3332
rect 31612 3278 31838 3330
rect 31890 3278 31892 3330
rect 31612 3276 31892 3278
rect 31612 800 31668 3276
rect 31836 3266 31892 3276
rect 32284 3330 32564 3332
rect 32284 3278 32510 3330
rect 32562 3278 32564 3330
rect 32284 3276 32564 3278
rect 32284 800 32340 3276
rect 32508 3266 32564 3276
rect 32956 3330 33236 3332
rect 32956 3278 33182 3330
rect 33234 3278 33236 3330
rect 32956 3276 33236 3278
rect 32956 800 33012 3276
rect 33180 3266 33236 3276
rect 33628 3330 33908 3332
rect 33628 3278 33854 3330
rect 33906 3278 33908 3330
rect 33628 3276 33908 3278
rect 33628 800 33684 3276
rect 33852 3266 33908 3276
rect 34300 3330 34580 3332
rect 34300 3278 34526 3330
rect 34578 3278 34580 3330
rect 34300 3276 34580 3278
rect 34300 800 34356 3276
rect 34524 3266 34580 3276
rect 34972 3330 35252 3332
rect 34972 3278 35198 3330
rect 35250 3278 35252 3330
rect 34972 3276 35252 3278
rect 34972 800 35028 3276
rect 35196 3266 35252 3276
rect 35644 3330 35924 3332
rect 35644 3278 35870 3330
rect 35922 3278 35924 3330
rect 35644 3276 35924 3278
rect 35644 800 35700 3276
rect 35868 3266 35924 3276
rect 36316 3330 36596 3332
rect 36316 3278 36542 3330
rect 36594 3278 36596 3330
rect 36316 3276 36596 3278
rect 36316 800 36372 3276
rect 36540 3266 36596 3276
rect 36988 3330 37268 3332
rect 36988 3278 37214 3330
rect 37266 3278 37268 3330
rect 36988 3276 37268 3278
rect 36988 800 37044 3276
rect 37212 3266 37268 3276
rect 37660 3330 37940 3332
rect 37660 3278 37886 3330
rect 37938 3278 37940 3330
rect 37660 3276 37940 3278
rect 37660 800 37716 3276
rect 37884 3266 37940 3276
rect 38332 3330 38612 3332
rect 38332 3278 38558 3330
rect 38610 3278 38612 3330
rect 38332 3276 38612 3278
rect 38332 800 38388 3276
rect 38556 3266 38612 3276
rect 39004 3330 39284 3332
rect 39004 3278 39230 3330
rect 39282 3278 39284 3330
rect 39004 3276 39284 3278
rect 39004 800 39060 3276
rect 39228 3266 39284 3276
rect 39676 3330 39956 3332
rect 39676 3278 39902 3330
rect 39954 3278 39956 3330
rect 39676 3276 39956 3278
rect 39676 800 39732 3276
rect 39900 3266 39956 3276
rect 40348 3330 40628 3332
rect 40348 3278 40574 3330
rect 40626 3278 40628 3330
rect 40348 3276 40628 3278
rect 40348 800 40404 3276
rect 40572 3266 40628 3276
rect 41692 3330 41748 3342
rect 41692 3278 41694 3330
rect 41746 3278 41748 3330
rect 41020 1762 41076 1774
rect 41020 1710 41022 1762
rect 41074 1710 41076 1762
rect 41020 800 41076 1710
rect 41692 1762 41748 3278
rect 41692 1710 41694 1762
rect 41746 1710 41748 1762
rect 41692 1698 41748 1710
rect 41804 3332 41860 3342
rect 41804 1540 41860 3276
rect 42364 3332 42420 3342
rect 42364 3238 42420 3276
rect 43036 3330 43092 3342
rect 43036 3278 43038 3330
rect 43090 3278 43092 3330
rect 41692 1484 41860 1540
rect 42364 1874 42420 1886
rect 42364 1822 42366 1874
rect 42418 1822 42420 1874
rect 41692 800 41748 1484
rect 42364 800 42420 1822
rect 43036 1874 43092 3278
rect 43036 1822 43038 1874
rect 43090 1822 43092 1874
rect 43036 1810 43092 1822
rect 43148 3332 43204 3342
rect 43148 1652 43204 3276
rect 43708 3332 43764 3342
rect 43708 3238 43764 3276
rect 44380 3330 44436 3342
rect 44380 3278 44382 3330
rect 44434 3278 44436 3330
rect 43036 1596 43204 1652
rect 43708 1762 43764 1774
rect 43708 1710 43710 1762
rect 43762 1710 43764 1762
rect 43036 800 43092 1596
rect 43708 800 43764 1710
rect 44380 1762 44436 3278
rect 45052 3330 45108 3342
rect 45052 3278 45054 3330
rect 45106 3278 45108 3330
rect 44380 1710 44382 1762
rect 44434 1710 44436 1762
rect 44380 1698 44436 1710
rect 44492 1874 44548 1886
rect 44492 1822 44494 1874
rect 44546 1822 44548 1874
rect 44492 1540 44548 1822
rect 45052 1874 45108 3278
rect 45052 1822 45054 1874
rect 45106 1822 45108 1874
rect 45052 1810 45108 1822
rect 45164 3332 45220 3342
rect 45164 1540 45220 3276
rect 45724 3332 45780 3342
rect 45724 3238 45780 3276
rect 46396 3330 46452 3342
rect 46396 3278 46398 3330
rect 46450 3278 46452 3330
rect 44380 1484 44548 1540
rect 45052 1484 45220 1540
rect 45724 1762 45780 1774
rect 45724 1710 45726 1762
rect 45778 1710 45780 1762
rect 44380 800 44436 1484
rect 45052 800 45108 1484
rect 45724 800 45780 1710
rect 46396 1762 46452 3278
rect 46396 1710 46398 1762
rect 46450 1710 46452 1762
rect 46396 1698 46452 1710
rect 46508 3332 46564 3342
rect 46508 1540 46564 3276
rect 47068 3332 47124 3342
rect 47068 3238 47124 3276
rect 47740 3330 47796 3342
rect 47740 3278 47742 3330
rect 47794 3278 47796 3330
rect 46396 1484 46564 1540
rect 47068 1762 47124 1774
rect 47068 1710 47070 1762
rect 47122 1710 47124 1762
rect 46396 800 46452 1484
rect 47068 800 47124 1710
rect 47740 1762 47796 3278
rect 48412 3330 48468 3342
rect 48412 3278 48414 3330
rect 48466 3278 48468 3330
rect 47740 1710 47742 1762
rect 47794 1710 47796 1762
rect 47740 1698 47796 1710
rect 47852 1874 47908 1886
rect 47852 1822 47854 1874
rect 47906 1822 47908 1874
rect 47852 1540 47908 1822
rect 48412 1874 48468 3278
rect 48412 1822 48414 1874
rect 48466 1822 48468 1874
rect 48412 1810 48468 1822
rect 48524 3332 48580 3342
rect 48524 1540 48580 3276
rect 49084 3332 49140 3342
rect 49084 3238 49140 3276
rect 49756 3330 49812 3342
rect 49756 3278 49758 3330
rect 49810 3278 49812 3330
rect 47740 1484 47908 1540
rect 48412 1484 48580 1540
rect 49084 1762 49140 1774
rect 49084 1710 49086 1762
rect 49138 1710 49140 1762
rect 47740 800 47796 1484
rect 48412 800 48468 1484
rect 49084 800 49140 1710
rect 49756 1762 49812 3278
rect 49756 1710 49758 1762
rect 49810 1710 49812 1762
rect 49756 1698 49812 1710
rect 49868 3332 49924 3342
rect 49868 1540 49924 3276
rect 50428 3332 50484 3342
rect 50428 3238 50484 3276
rect 51100 3330 51156 3342
rect 51100 3278 51102 3330
rect 51154 3278 51156 3330
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 49756 1484 49924 1540
rect 50428 1762 50484 1774
rect 50428 1710 50430 1762
rect 50482 1710 50484 1762
rect 49756 800 49812 1484
rect 50428 800 50484 1710
rect 51100 1762 51156 3278
rect 51772 3330 51828 3342
rect 51772 3278 51774 3330
rect 51826 3278 51828 3330
rect 51100 1710 51102 1762
rect 51154 1710 51156 1762
rect 51100 1698 51156 1710
rect 51212 1874 51268 1886
rect 51212 1822 51214 1874
rect 51266 1822 51268 1874
rect 51212 1540 51268 1822
rect 51772 1874 51828 3278
rect 51772 1822 51774 1874
rect 51826 1822 51828 1874
rect 51772 1810 51828 1822
rect 51884 3332 51940 3342
rect 51884 1540 51940 3276
rect 52444 3332 52500 3342
rect 52444 3238 52500 3276
rect 53116 3330 53172 3342
rect 53116 3278 53118 3330
rect 53170 3278 53172 3330
rect 51100 1484 51268 1540
rect 51772 1484 51940 1540
rect 52444 1762 52500 1774
rect 52444 1710 52446 1762
rect 52498 1710 52500 1762
rect 51100 800 51156 1484
rect 51772 800 51828 1484
rect 52444 800 52500 1710
rect 53116 1762 53172 3278
rect 53116 1710 53118 1762
rect 53170 1710 53172 1762
rect 53116 1698 53172 1710
rect 53228 3332 53284 3342
rect 53228 1540 53284 3276
rect 53788 3332 53844 3342
rect 53788 3238 53844 3276
rect 54460 3330 54516 3342
rect 54460 3278 54462 3330
rect 54514 3278 54516 3330
rect 53116 1484 53284 1540
rect 53788 1762 53844 1774
rect 53788 1710 53790 1762
rect 53842 1710 53844 1762
rect 53116 800 53172 1484
rect 53788 800 53844 1710
rect 54460 1762 54516 3278
rect 55132 3330 55188 3342
rect 55132 3278 55134 3330
rect 55186 3278 55188 3330
rect 54460 1710 54462 1762
rect 54514 1710 54516 1762
rect 54460 1698 54516 1710
rect 54572 1986 54628 1998
rect 54572 1934 54574 1986
rect 54626 1934 54628 1986
rect 54572 1540 54628 1934
rect 55132 1986 55188 3278
rect 55132 1934 55134 1986
rect 55186 1934 55188 1986
rect 55132 1922 55188 1934
rect 55804 3330 55860 3342
rect 55804 3278 55806 3330
rect 55858 3278 55860 3330
rect 54460 1484 54628 1540
rect 55132 1764 55188 1774
rect 54460 800 54516 1484
rect 55132 800 55188 1708
rect 55804 1764 55860 3278
rect 56476 3330 56532 3342
rect 56476 3278 56478 3330
rect 56530 3278 56532 3330
rect 55804 1698 55860 1708
rect 55916 1762 55972 1774
rect 55916 1710 55918 1762
rect 55970 1710 55972 1762
rect 55916 1540 55972 1710
rect 56476 1762 56532 3278
rect 56476 1710 56478 1762
rect 56530 1710 56532 1762
rect 56476 1698 56532 1710
rect 56588 3332 56644 3342
rect 56588 1540 56644 3276
rect 57148 3332 57204 3342
rect 57148 3238 57204 3276
rect 57820 3330 57876 3342
rect 57820 3278 57822 3330
rect 57874 3278 57876 3330
rect 55804 1484 55972 1540
rect 56476 1484 56644 1540
rect 57148 1762 57204 1774
rect 57148 1710 57150 1762
rect 57202 1710 57204 1762
rect 55804 800 55860 1484
rect 56476 800 56532 1484
rect 57148 800 57204 1710
rect 57820 1762 57876 3278
rect 58492 3330 58548 3342
rect 58492 3278 58494 3330
rect 58546 3278 58548 3330
rect 57820 1710 57822 1762
rect 57874 1710 57876 1762
rect 57820 1698 57876 1710
rect 57932 1874 57988 1886
rect 57932 1822 57934 1874
rect 57986 1822 57988 1874
rect 57932 1540 57988 1822
rect 58492 1874 58548 3278
rect 58492 1822 58494 1874
rect 58546 1822 58548 1874
rect 58492 1810 58548 1822
rect 58604 3332 58660 3342
rect 58604 1540 58660 3276
rect 59164 3332 59220 3342
rect 59164 3238 59220 3276
rect 59836 3330 59892 3342
rect 59836 3278 59838 3330
rect 59890 3278 59892 3330
rect 57820 1484 57988 1540
rect 58492 1484 58660 1540
rect 59164 1762 59220 1774
rect 59164 1710 59166 1762
rect 59218 1710 59220 1762
rect 57820 800 57876 1484
rect 58492 800 58548 1484
rect 59164 800 59220 1710
rect 59836 1762 59892 3278
rect 59836 1710 59838 1762
rect 59890 1710 59892 1762
rect 59836 1698 59892 1710
rect 59948 3332 60004 3342
rect 59948 1540 60004 3276
rect 60508 3332 60564 3342
rect 60508 3238 60564 3276
rect 61180 3332 61236 3342
rect 59836 1484 60004 1540
rect 60508 1762 60564 1774
rect 60508 1710 60510 1762
rect 60562 1710 60564 1762
rect 59836 800 59892 1484
rect 60508 800 60564 1710
rect 61180 800 61236 3276
rect 61628 3330 61684 3342
rect 61628 3278 61630 3330
rect 61682 3278 61684 3330
rect 61628 1762 61684 3278
rect 62300 3332 62356 3342
rect 62300 3238 62356 3276
rect 62972 3330 63028 3342
rect 62972 3278 62974 3330
rect 63026 3278 63028 3330
rect 61628 1710 61630 1762
rect 61682 1710 61684 1762
rect 61628 1698 61684 1710
rect 61852 1764 61908 1774
rect 61852 800 61908 1708
rect 62524 1762 62580 1774
rect 62524 1710 62526 1762
rect 62578 1710 62580 1762
rect 62524 800 62580 1710
rect 62972 1764 63028 3278
rect 62972 1698 63028 1708
rect 63196 3332 63252 3342
rect 63196 800 63252 3276
rect 63644 3330 63700 3342
rect 63644 3278 63646 3330
rect 63698 3278 63700 3330
rect 63644 1762 63700 3278
rect 64316 3332 64372 3342
rect 64316 3238 64372 3276
rect 64540 3332 64596 3342
rect 63644 1710 63646 1762
rect 63698 1710 63700 1762
rect 63644 1698 63700 1710
rect 63868 1762 63924 1774
rect 63868 1710 63870 1762
rect 63922 1710 63924 1762
rect 63868 800 63924 1710
rect 64540 800 64596 3276
rect 64988 3330 65044 3342
rect 64988 3278 64990 3330
rect 65042 3278 65044 3330
rect 64988 1762 65044 3278
rect 65660 3332 65716 3342
rect 65660 3238 65716 3276
rect 66332 3330 66388 3342
rect 66332 3278 66334 3330
rect 66386 3278 66388 3330
rect 64988 1710 64990 1762
rect 65042 1710 65044 1762
rect 64988 1698 65044 1710
rect 65212 1764 65268 1774
rect 65212 800 65268 1708
rect 65884 1762 65940 1774
rect 65884 1710 65886 1762
rect 65938 1710 65940 1762
rect 65884 800 65940 1710
rect 66332 1764 66388 3278
rect 66332 1698 66388 1708
rect 66556 3332 66612 3342
rect 66556 800 66612 3276
rect 67004 3330 67060 3342
rect 67004 3278 67006 3330
rect 67058 3278 67060 3330
rect 67004 1762 67060 3278
rect 67676 3332 67732 3342
rect 67676 3238 67732 3276
rect 67900 3332 67956 3342
rect 67004 1710 67006 1762
rect 67058 1710 67060 1762
rect 67004 1698 67060 1710
rect 67228 1762 67284 1774
rect 67228 1710 67230 1762
rect 67282 1710 67284 1762
rect 67228 800 67284 1710
rect 67900 800 67956 3276
rect 68348 3330 68404 3342
rect 68348 3278 68350 3330
rect 68402 3278 68404 3330
rect 68348 1762 68404 3278
rect 69020 3332 69076 3342
rect 69020 3238 69076 3276
rect 69692 3330 69748 3342
rect 69692 3278 69694 3330
rect 69746 3278 69748 3330
rect 68348 1710 68350 1762
rect 68402 1710 68404 1762
rect 68348 1698 68404 1710
rect 68572 1764 68628 1774
rect 68572 800 68628 1708
rect 69244 1762 69300 1774
rect 69244 1710 69246 1762
rect 69298 1710 69300 1762
rect 69244 800 69300 1710
rect 69692 1764 69748 3278
rect 69692 1698 69748 1708
rect 69916 3332 69972 3342
rect 69916 800 69972 3276
rect 70364 3330 70420 3342
rect 70364 3278 70366 3330
rect 70418 3278 70420 3330
rect 70364 1762 70420 3278
rect 71036 3332 71092 3342
rect 71036 3238 71092 3276
rect 71260 3332 71316 3342
rect 70364 1710 70366 1762
rect 70418 1710 70420 1762
rect 70364 1698 70420 1710
rect 70588 1762 70644 1774
rect 70588 1710 70590 1762
rect 70642 1710 70644 1762
rect 70588 800 70644 1710
rect 71260 800 71316 3276
rect 71708 3330 71764 3342
rect 71708 3278 71710 3330
rect 71762 3278 71764 3330
rect 71708 1762 71764 3278
rect 72380 3332 72436 3342
rect 72380 3238 72436 3276
rect 73052 3330 73108 3342
rect 73052 3278 73054 3330
rect 73106 3278 73108 3330
rect 71708 1710 71710 1762
rect 71762 1710 71764 1762
rect 71708 1698 71764 1710
rect 71932 1764 71988 1774
rect 71932 800 71988 1708
rect 72604 1762 72660 1774
rect 72604 1710 72606 1762
rect 72658 1710 72660 1762
rect 72604 800 72660 1710
rect 73052 1764 73108 3278
rect 73052 1698 73108 1708
rect 73164 1540 73220 4396
rect 73276 4386 73332 4396
rect 73500 4450 74004 4452
rect 73500 4398 73950 4450
rect 74002 4398 74004 4450
rect 73500 4396 74004 4398
rect 73052 1484 73220 1540
rect 73388 3332 73444 3342
rect 73052 800 73108 1484
rect 73388 980 73444 3276
rect 73276 924 73444 980
rect 73276 800 73332 924
rect 73500 800 73556 4396
rect 73948 4386 74004 4396
rect 73724 3330 73780 3342
rect 73724 3278 73726 3330
rect 73778 3278 73780 3330
rect 73724 1762 73780 3278
rect 74396 3332 74452 3342
rect 74396 3238 74452 3276
rect 73724 1710 73726 1762
rect 73778 1710 73780 1762
rect 73724 1698 73780 1710
rect 6272 0 6384 800
rect 6496 0 6608 800
rect 6720 0 6832 800
rect 6944 0 7056 800
rect 7168 0 7280 800
rect 7392 0 7504 800
rect 7616 0 7728 800
rect 7840 0 7952 800
rect 8064 0 8176 800
rect 8288 0 8400 800
rect 8512 0 8624 800
rect 8736 0 8848 800
rect 8960 0 9072 800
rect 9184 0 9296 800
rect 9408 0 9520 800
rect 9632 0 9744 800
rect 9856 0 9968 800
rect 10080 0 10192 800
rect 10304 0 10416 800
rect 10528 0 10640 800
rect 10752 0 10864 800
rect 10976 0 11088 800
rect 11200 0 11312 800
rect 11424 0 11536 800
rect 11648 0 11760 800
rect 11872 0 11984 800
rect 12096 0 12208 800
rect 12320 0 12432 800
rect 12544 0 12656 800
rect 12768 0 12880 800
rect 12992 0 13104 800
rect 13216 0 13328 800
rect 13440 0 13552 800
rect 13664 0 13776 800
rect 13888 0 14000 800
rect 14112 0 14224 800
rect 14336 0 14448 800
rect 14560 0 14672 800
rect 14784 0 14896 800
rect 15008 0 15120 800
rect 15232 0 15344 800
rect 15456 0 15568 800
rect 15680 0 15792 800
rect 15904 0 16016 800
rect 16128 0 16240 800
rect 16352 0 16464 800
rect 16576 0 16688 800
rect 16800 0 16912 800
rect 17024 0 17136 800
rect 17248 0 17360 800
rect 17472 0 17584 800
rect 17696 0 17808 800
rect 17920 0 18032 800
rect 18144 0 18256 800
rect 18368 0 18480 800
rect 18592 0 18704 800
rect 18816 0 18928 800
rect 19040 0 19152 800
rect 19264 0 19376 800
rect 19488 0 19600 800
rect 19712 0 19824 800
rect 19936 0 20048 800
rect 20160 0 20272 800
rect 20384 0 20496 800
rect 20608 0 20720 800
rect 20832 0 20944 800
rect 21056 0 21168 800
rect 21280 0 21392 800
rect 21504 0 21616 800
rect 21728 0 21840 800
rect 21952 0 22064 800
rect 22176 0 22288 800
rect 22400 0 22512 800
rect 22624 0 22736 800
rect 22848 0 22960 800
rect 23072 0 23184 800
rect 23296 0 23408 800
rect 23520 0 23632 800
rect 23744 0 23856 800
rect 23968 0 24080 800
rect 24192 0 24304 800
rect 24416 0 24528 800
rect 24640 0 24752 800
rect 24864 0 24976 800
rect 25088 0 25200 800
rect 25312 0 25424 800
rect 25536 0 25648 800
rect 25760 0 25872 800
rect 25984 0 26096 800
rect 26208 0 26320 800
rect 26432 0 26544 800
rect 26656 0 26768 800
rect 26880 0 26992 800
rect 27104 0 27216 800
rect 27328 0 27440 800
rect 27552 0 27664 800
rect 27776 0 27888 800
rect 28000 0 28112 800
rect 28224 0 28336 800
rect 28448 0 28560 800
rect 28672 0 28784 800
rect 28896 0 29008 800
rect 29120 0 29232 800
rect 29344 0 29456 800
rect 29568 0 29680 800
rect 29792 0 29904 800
rect 30016 0 30128 800
rect 30240 0 30352 800
rect 30464 0 30576 800
rect 30688 0 30800 800
rect 30912 0 31024 800
rect 31136 0 31248 800
rect 31360 0 31472 800
rect 31584 0 31696 800
rect 31808 0 31920 800
rect 32032 0 32144 800
rect 32256 0 32368 800
rect 32480 0 32592 800
rect 32704 0 32816 800
rect 32928 0 33040 800
rect 33152 0 33264 800
rect 33376 0 33488 800
rect 33600 0 33712 800
rect 33824 0 33936 800
rect 34048 0 34160 800
rect 34272 0 34384 800
rect 34496 0 34608 800
rect 34720 0 34832 800
rect 34944 0 35056 800
rect 35168 0 35280 800
rect 35392 0 35504 800
rect 35616 0 35728 800
rect 35840 0 35952 800
rect 36064 0 36176 800
rect 36288 0 36400 800
rect 36512 0 36624 800
rect 36736 0 36848 800
rect 36960 0 37072 800
rect 37184 0 37296 800
rect 37408 0 37520 800
rect 37632 0 37744 800
rect 37856 0 37968 800
rect 38080 0 38192 800
rect 38304 0 38416 800
rect 38528 0 38640 800
rect 38752 0 38864 800
rect 38976 0 39088 800
rect 39200 0 39312 800
rect 39424 0 39536 800
rect 39648 0 39760 800
rect 39872 0 39984 800
rect 40096 0 40208 800
rect 40320 0 40432 800
rect 40544 0 40656 800
rect 40768 0 40880 800
rect 40992 0 41104 800
rect 41216 0 41328 800
rect 41440 0 41552 800
rect 41664 0 41776 800
rect 41888 0 42000 800
rect 42112 0 42224 800
rect 42336 0 42448 800
rect 42560 0 42672 800
rect 42784 0 42896 800
rect 43008 0 43120 800
rect 43232 0 43344 800
rect 43456 0 43568 800
rect 43680 0 43792 800
rect 43904 0 44016 800
rect 44128 0 44240 800
rect 44352 0 44464 800
rect 44576 0 44688 800
rect 44800 0 44912 800
rect 45024 0 45136 800
rect 45248 0 45360 800
rect 45472 0 45584 800
rect 45696 0 45808 800
rect 45920 0 46032 800
rect 46144 0 46256 800
rect 46368 0 46480 800
rect 46592 0 46704 800
rect 46816 0 46928 800
rect 47040 0 47152 800
rect 47264 0 47376 800
rect 47488 0 47600 800
rect 47712 0 47824 800
rect 47936 0 48048 800
rect 48160 0 48272 800
rect 48384 0 48496 800
rect 48608 0 48720 800
rect 48832 0 48944 800
rect 49056 0 49168 800
rect 49280 0 49392 800
rect 49504 0 49616 800
rect 49728 0 49840 800
rect 49952 0 50064 800
rect 50176 0 50288 800
rect 50400 0 50512 800
rect 50624 0 50736 800
rect 50848 0 50960 800
rect 51072 0 51184 800
rect 51296 0 51408 800
rect 51520 0 51632 800
rect 51744 0 51856 800
rect 51968 0 52080 800
rect 52192 0 52304 800
rect 52416 0 52528 800
rect 52640 0 52752 800
rect 52864 0 52976 800
rect 53088 0 53200 800
rect 53312 0 53424 800
rect 53536 0 53648 800
rect 53760 0 53872 800
rect 53984 0 54096 800
rect 54208 0 54320 800
rect 54432 0 54544 800
rect 54656 0 54768 800
rect 54880 0 54992 800
rect 55104 0 55216 800
rect 55328 0 55440 800
rect 55552 0 55664 800
rect 55776 0 55888 800
rect 56000 0 56112 800
rect 56224 0 56336 800
rect 56448 0 56560 800
rect 56672 0 56784 800
rect 56896 0 57008 800
rect 57120 0 57232 800
rect 57344 0 57456 800
rect 57568 0 57680 800
rect 57792 0 57904 800
rect 58016 0 58128 800
rect 58240 0 58352 800
rect 58464 0 58576 800
rect 58688 0 58800 800
rect 58912 0 59024 800
rect 59136 0 59248 800
rect 59360 0 59472 800
rect 59584 0 59696 800
rect 59808 0 59920 800
rect 60032 0 60144 800
rect 60256 0 60368 800
rect 60480 0 60592 800
rect 60704 0 60816 800
rect 60928 0 61040 800
rect 61152 0 61264 800
rect 61376 0 61488 800
rect 61600 0 61712 800
rect 61824 0 61936 800
rect 62048 0 62160 800
rect 62272 0 62384 800
rect 62496 0 62608 800
rect 62720 0 62832 800
rect 62944 0 63056 800
rect 63168 0 63280 800
rect 63392 0 63504 800
rect 63616 0 63728 800
rect 63840 0 63952 800
rect 64064 0 64176 800
rect 64288 0 64400 800
rect 64512 0 64624 800
rect 64736 0 64848 800
rect 64960 0 65072 800
rect 65184 0 65296 800
rect 65408 0 65520 800
rect 65632 0 65744 800
rect 65856 0 65968 800
rect 66080 0 66192 800
rect 66304 0 66416 800
rect 66528 0 66640 800
rect 66752 0 66864 800
rect 66976 0 67088 800
rect 67200 0 67312 800
rect 67424 0 67536 800
rect 67648 0 67760 800
rect 67872 0 67984 800
rect 68096 0 68208 800
rect 68320 0 68432 800
rect 68544 0 68656 800
rect 68768 0 68880 800
rect 68992 0 69104 800
rect 69216 0 69328 800
rect 69440 0 69552 800
rect 69664 0 69776 800
rect 69888 0 70000 800
rect 70112 0 70224 800
rect 70336 0 70448 800
rect 70560 0 70672 800
rect 70784 0 70896 800
rect 71008 0 71120 800
rect 71232 0 71344 800
rect 71456 0 71568 800
rect 71680 0 71792 800
rect 71904 0 72016 800
rect 72128 0 72240 800
rect 72352 0 72464 800
rect 72576 0 72688 800
rect 72800 0 72912 800
rect 73024 0 73136 800
rect 73248 0 73360 800
rect 73472 0 73584 800
<< via2 >>
rect 4476 76074 4532 76076
rect 4476 76022 4478 76074
rect 4478 76022 4530 76074
rect 4530 76022 4532 76074
rect 4476 76020 4532 76022
rect 4580 76074 4636 76076
rect 4580 76022 4582 76074
rect 4582 76022 4634 76074
rect 4634 76022 4636 76074
rect 4580 76020 4636 76022
rect 4684 76074 4740 76076
rect 4684 76022 4686 76074
rect 4686 76022 4738 76074
rect 4738 76022 4740 76074
rect 4684 76020 4740 76022
rect 3388 75852 3444 75908
rect 6524 77308 6580 77364
rect 5068 76466 5124 76468
rect 5068 76414 5070 76466
rect 5070 76414 5122 76466
rect 5122 76414 5124 76466
rect 5068 76412 5124 76414
rect 6524 76412 6580 76468
rect 13132 76466 13188 76468
rect 13132 76414 13134 76466
rect 13134 76414 13186 76466
rect 13186 76414 13188 76466
rect 13132 76412 13188 76414
rect 13804 76412 13860 76468
rect 4476 74506 4532 74508
rect 4476 74454 4478 74506
rect 4478 74454 4530 74506
rect 4530 74454 4532 74506
rect 4476 74452 4532 74454
rect 4580 74506 4636 74508
rect 4580 74454 4582 74506
rect 4582 74454 4634 74506
rect 4634 74454 4636 74506
rect 4580 74452 4636 74454
rect 4684 74506 4740 74508
rect 4684 74454 4686 74506
rect 4686 74454 4738 74506
rect 4738 74454 4740 74506
rect 4684 74452 4740 74454
rect 4476 72938 4532 72940
rect 4476 72886 4478 72938
rect 4478 72886 4530 72938
rect 4530 72886 4532 72938
rect 4476 72884 4532 72886
rect 4580 72938 4636 72940
rect 4580 72886 4582 72938
rect 4582 72886 4634 72938
rect 4634 72886 4636 72938
rect 4580 72884 4636 72886
rect 4684 72938 4740 72940
rect 4684 72886 4686 72938
rect 4686 72886 4738 72938
rect 4738 72886 4740 72938
rect 4684 72884 4740 72886
rect 15148 76466 15204 76468
rect 15148 76414 15150 76466
rect 15150 76414 15202 76466
rect 15202 76414 15204 76466
rect 15148 76412 15204 76414
rect 15820 76412 15876 76468
rect 16940 75628 16996 75684
rect 17836 75682 17892 75684
rect 17836 75630 17838 75682
rect 17838 75630 17890 75682
rect 17890 75630 17892 75682
rect 17836 75628 17892 75630
rect 19836 76858 19892 76860
rect 19836 76806 19838 76858
rect 19838 76806 19890 76858
rect 19890 76806 19892 76858
rect 19836 76804 19892 76806
rect 19940 76858 19996 76860
rect 19940 76806 19942 76858
rect 19942 76806 19994 76858
rect 19994 76806 19996 76858
rect 19940 76804 19996 76806
rect 20044 76858 20100 76860
rect 20044 76806 20046 76858
rect 20046 76806 20098 76858
rect 20098 76806 20100 76858
rect 20044 76804 20100 76806
rect 20972 76188 21028 76244
rect 19180 75740 19236 75796
rect 19852 75794 19908 75796
rect 19852 75742 19854 75794
rect 19854 75742 19906 75794
rect 19906 75742 19908 75794
rect 19852 75740 19908 75742
rect 19836 75290 19892 75292
rect 19836 75238 19838 75290
rect 19838 75238 19890 75290
rect 19890 75238 19892 75290
rect 19836 75236 19892 75238
rect 19940 75290 19996 75292
rect 19940 75238 19942 75290
rect 19942 75238 19994 75290
rect 19994 75238 19996 75290
rect 19940 75236 19996 75238
rect 20044 75290 20100 75292
rect 20044 75238 20046 75290
rect 20046 75238 20098 75290
rect 20098 75238 20100 75290
rect 20044 75236 20100 75238
rect 21084 75516 21140 75572
rect 21644 75852 21700 75908
rect 20188 75068 20244 75124
rect 21756 75570 21812 75572
rect 21756 75518 21758 75570
rect 21758 75518 21810 75570
rect 21810 75518 21812 75570
rect 21756 75516 21812 75518
rect 25004 76466 25060 76468
rect 25004 76414 25006 76466
rect 25006 76414 25058 76466
rect 25058 76414 25060 76466
rect 25004 76412 25060 76414
rect 23212 76076 23268 76132
rect 23996 76076 24052 76132
rect 26796 76524 26852 76580
rect 27244 76524 27300 76580
rect 27804 76300 27860 76356
rect 21644 74956 21700 75012
rect 29260 76412 29316 76468
rect 28812 76354 28868 76356
rect 28812 76302 28814 76354
rect 28814 76302 28866 76354
rect 28866 76302 28868 76354
rect 28812 76300 28868 76302
rect 29820 76300 29876 76356
rect 29484 75964 29540 76020
rect 29372 75794 29428 75796
rect 29372 75742 29374 75794
rect 29374 75742 29426 75794
rect 29426 75742 29428 75794
rect 29372 75740 29428 75742
rect 28588 74284 28644 74340
rect 28924 74732 28980 74788
rect 30716 76354 30772 76356
rect 30716 76302 30718 76354
rect 30718 76302 30770 76354
rect 30770 76302 30772 76354
rect 30716 76300 30772 76302
rect 33180 77532 33236 77588
rect 33068 76524 33124 76580
rect 31836 76300 31892 76356
rect 30828 75740 30884 75796
rect 30044 75682 30100 75684
rect 30044 75630 30046 75682
rect 30046 75630 30098 75682
rect 30098 75630 30100 75682
rect 30044 75628 30100 75630
rect 30268 75516 30324 75572
rect 29932 75010 29988 75012
rect 29932 74958 29934 75010
rect 29934 74958 29986 75010
rect 29986 74958 29988 75010
rect 29932 74956 29988 74958
rect 29372 74844 29428 74900
rect 29260 74786 29316 74788
rect 29260 74734 29262 74786
rect 29262 74734 29314 74786
rect 29314 74734 29316 74786
rect 29260 74732 29316 74734
rect 29820 74226 29876 74228
rect 29820 74174 29822 74226
rect 29822 74174 29874 74226
rect 29874 74174 29876 74226
rect 29820 74172 29876 74174
rect 29148 73836 29204 73892
rect 30268 73890 30324 73892
rect 30268 73838 30270 73890
rect 30270 73838 30322 73890
rect 30322 73838 30324 73890
rect 30268 73836 30324 73838
rect 19836 73722 19892 73724
rect 19836 73670 19838 73722
rect 19838 73670 19890 73722
rect 19890 73670 19892 73722
rect 19836 73668 19892 73670
rect 19940 73722 19996 73724
rect 19940 73670 19942 73722
rect 19942 73670 19994 73722
rect 19994 73670 19996 73722
rect 19940 73668 19996 73670
rect 20044 73722 20100 73724
rect 20044 73670 20046 73722
rect 20046 73670 20098 73722
rect 20098 73670 20100 73722
rect 20044 73668 20100 73670
rect 30492 75628 30548 75684
rect 30604 75516 30660 75572
rect 31164 75516 31220 75572
rect 31276 75404 31332 75460
rect 31388 75180 31444 75236
rect 31164 74956 31220 75012
rect 31052 74172 31108 74228
rect 30380 72604 30436 72660
rect 32732 76354 32788 76356
rect 32732 76302 32734 76354
rect 32734 76302 32786 76354
rect 32786 76302 32788 76354
rect 32732 76300 32788 76302
rect 32172 75964 32228 76020
rect 31836 75180 31892 75236
rect 31836 74172 31892 74228
rect 32060 75516 32116 75572
rect 32620 75570 32676 75572
rect 32620 75518 32622 75570
rect 32622 75518 32674 75570
rect 32674 75518 32676 75570
rect 32620 75516 32676 75518
rect 32060 74898 32116 74900
rect 32060 74846 32062 74898
rect 32062 74846 32114 74898
rect 32114 74846 32116 74898
rect 32060 74844 32116 74846
rect 32284 74786 32340 74788
rect 32284 74734 32286 74786
rect 32286 74734 32338 74786
rect 32338 74734 32340 74786
rect 32284 74732 32340 74734
rect 31500 73890 31556 73892
rect 31500 73838 31502 73890
rect 31502 73838 31554 73890
rect 31554 73838 31556 73890
rect 31500 73836 31556 73838
rect 32508 75180 32564 75236
rect 33180 75404 33236 75460
rect 33180 75180 33236 75236
rect 33292 75068 33348 75124
rect 32732 74060 32788 74116
rect 33516 74674 33572 74676
rect 33516 74622 33518 74674
rect 33518 74622 33570 74674
rect 33570 74622 33572 74674
rect 33516 74620 33572 74622
rect 33852 75516 33908 75572
rect 33740 74898 33796 74900
rect 33740 74846 33742 74898
rect 33742 74846 33794 74898
rect 33794 74846 33796 74898
rect 33740 74844 33796 74846
rect 33404 74060 33460 74116
rect 31276 72604 31332 72660
rect 31836 72604 31892 72660
rect 15820 72268 15876 72324
rect 19836 72154 19892 72156
rect 19836 72102 19838 72154
rect 19838 72102 19890 72154
rect 19890 72102 19892 72154
rect 19836 72100 19892 72102
rect 19940 72154 19996 72156
rect 19940 72102 19942 72154
rect 19942 72102 19994 72154
rect 19994 72102 19996 72154
rect 19940 72100 19996 72102
rect 20044 72154 20100 72156
rect 20044 72102 20046 72154
rect 20046 72102 20098 72154
rect 20098 72102 20100 72154
rect 20044 72100 20100 72102
rect 13804 71484 13860 71540
rect 4476 71370 4532 71372
rect 4476 71318 4478 71370
rect 4478 71318 4530 71370
rect 4530 71318 4532 71370
rect 4476 71316 4532 71318
rect 4580 71370 4636 71372
rect 4580 71318 4582 71370
rect 4582 71318 4634 71370
rect 4634 71318 4636 71370
rect 4580 71316 4636 71318
rect 4684 71370 4740 71372
rect 4684 71318 4686 71370
rect 4686 71318 4738 71370
rect 4738 71318 4740 71370
rect 4684 71316 4740 71318
rect 19836 70586 19892 70588
rect 19836 70534 19838 70586
rect 19838 70534 19890 70586
rect 19890 70534 19892 70586
rect 19836 70532 19892 70534
rect 19940 70586 19996 70588
rect 19940 70534 19942 70586
rect 19942 70534 19994 70586
rect 19994 70534 19996 70586
rect 19940 70532 19996 70534
rect 20044 70586 20100 70588
rect 20044 70534 20046 70586
rect 20046 70534 20098 70586
rect 20098 70534 20100 70586
rect 20044 70532 20100 70534
rect 31948 72658 32004 72660
rect 31948 72606 31950 72658
rect 31950 72606 32002 72658
rect 32002 72606 32004 72658
rect 31948 72604 32004 72606
rect 34636 76412 34692 76468
rect 34076 75516 34132 75572
rect 34412 75570 34468 75572
rect 34412 75518 34414 75570
rect 34414 75518 34466 75570
rect 34466 75518 34468 75570
rect 34412 75516 34468 75518
rect 34300 75404 34356 75460
rect 33964 74338 34020 74340
rect 33964 74286 33966 74338
rect 33966 74286 34018 74338
rect 34018 74286 34020 74338
rect 33964 74284 34020 74286
rect 35756 77196 35812 77252
rect 34188 73724 34244 73780
rect 34412 74284 34468 74340
rect 34524 74226 34580 74228
rect 34524 74174 34526 74226
rect 34526 74174 34578 74226
rect 34578 74174 34580 74226
rect 34524 74172 34580 74174
rect 34188 72658 34244 72660
rect 34188 72606 34190 72658
rect 34190 72606 34242 72658
rect 34242 72606 34244 72658
rect 34188 72604 34244 72606
rect 35084 76188 35140 76244
rect 35196 76074 35252 76076
rect 35196 76022 35198 76074
rect 35198 76022 35250 76074
rect 35250 76022 35252 76074
rect 35196 76020 35252 76022
rect 35300 76074 35356 76076
rect 35300 76022 35302 76074
rect 35302 76022 35354 76074
rect 35354 76022 35356 76074
rect 35300 76020 35356 76022
rect 35404 76074 35460 76076
rect 35404 76022 35406 76074
rect 35406 76022 35458 76074
rect 35458 76022 35460 76074
rect 35404 76020 35460 76022
rect 34972 75404 35028 75460
rect 35196 74898 35252 74900
rect 35196 74846 35198 74898
rect 35198 74846 35250 74898
rect 35250 74846 35252 74898
rect 35196 74844 35252 74846
rect 36092 76466 36148 76468
rect 36092 76414 36094 76466
rect 36094 76414 36146 76466
rect 36146 76414 36148 76466
rect 36092 76412 36148 76414
rect 35756 75404 35812 75460
rect 35980 76188 36036 76244
rect 35532 74732 35588 74788
rect 35196 74506 35252 74508
rect 35196 74454 35198 74506
rect 35198 74454 35250 74506
rect 35250 74454 35252 74506
rect 35196 74452 35252 74454
rect 35300 74506 35356 74508
rect 35300 74454 35302 74506
rect 35302 74454 35354 74506
rect 35354 74454 35356 74506
rect 35300 74452 35356 74454
rect 35404 74506 35460 74508
rect 35404 74454 35406 74506
rect 35406 74454 35458 74506
rect 35458 74454 35460 74506
rect 35404 74452 35460 74454
rect 35084 74338 35140 74340
rect 35084 74286 35086 74338
rect 35086 74286 35138 74338
rect 35138 74286 35140 74338
rect 35084 74284 35140 74286
rect 35644 74844 35700 74900
rect 35644 74226 35700 74228
rect 35644 74174 35646 74226
rect 35646 74174 35698 74226
rect 35698 74174 35700 74226
rect 35644 74172 35700 74174
rect 35308 74060 35364 74116
rect 35756 74396 35812 74452
rect 36652 76076 36708 76132
rect 36316 75852 36372 75908
rect 35532 73052 35588 73108
rect 35196 72938 35252 72940
rect 35196 72886 35198 72938
rect 35198 72886 35250 72938
rect 35250 72886 35252 72938
rect 35196 72884 35252 72886
rect 35300 72938 35356 72940
rect 35300 72886 35302 72938
rect 35302 72886 35354 72938
rect 35354 72886 35356 72938
rect 35300 72884 35356 72886
rect 35404 72938 35460 72940
rect 35404 72886 35406 72938
rect 35406 72886 35458 72938
rect 35458 72886 35460 72938
rect 35404 72884 35460 72886
rect 35420 72658 35476 72660
rect 35420 72606 35422 72658
rect 35422 72606 35474 72658
rect 35474 72606 35476 72658
rect 35420 72604 35476 72606
rect 35308 72322 35364 72324
rect 35308 72270 35310 72322
rect 35310 72270 35362 72322
rect 35362 72270 35364 72322
rect 35308 72268 35364 72270
rect 34860 71538 34916 71540
rect 34860 71486 34862 71538
rect 34862 71486 34914 71538
rect 34914 71486 34916 71538
rect 34860 71484 34916 71486
rect 35196 71370 35252 71372
rect 35196 71318 35198 71370
rect 35198 71318 35250 71370
rect 35250 71318 35252 71370
rect 35196 71316 35252 71318
rect 35300 71370 35356 71372
rect 35300 71318 35302 71370
rect 35302 71318 35354 71370
rect 35354 71318 35356 71370
rect 35300 71316 35356 71318
rect 35404 71370 35460 71372
rect 35404 71318 35406 71370
rect 35406 71318 35458 71370
rect 35458 71318 35460 71370
rect 35404 71316 35460 71318
rect 34300 71036 34356 71092
rect 35196 71090 35252 71092
rect 35196 71038 35198 71090
rect 35198 71038 35250 71090
rect 35250 71038 35252 71090
rect 35196 71036 35252 71038
rect 35644 71090 35700 71092
rect 35644 71038 35646 71090
rect 35646 71038 35698 71090
rect 35698 71038 35700 71090
rect 35644 71036 35700 71038
rect 36092 70924 36148 70980
rect 36540 74956 36596 75012
rect 36316 74620 36372 74676
rect 36316 73948 36372 74004
rect 36428 72434 36484 72436
rect 36428 72382 36430 72434
rect 36430 72382 36482 72434
rect 36482 72382 36484 72434
rect 36428 72380 36484 72382
rect 36428 71986 36484 71988
rect 36428 71934 36430 71986
rect 36430 71934 36482 71986
rect 36482 71934 36484 71986
rect 36428 71932 36484 71934
rect 36204 71260 36260 71316
rect 36428 70978 36484 70980
rect 36428 70926 36430 70978
rect 36430 70926 36482 70978
rect 36482 70926 36484 70978
rect 36428 70924 36484 70926
rect 35532 70476 35588 70532
rect 31836 70364 31892 70420
rect 36876 74732 36932 74788
rect 37884 76748 37940 76804
rect 38332 76636 38388 76692
rect 37548 75458 37604 75460
rect 37548 75406 37550 75458
rect 37550 75406 37602 75458
rect 37602 75406 37604 75458
rect 37548 75404 37604 75406
rect 37548 75180 37604 75236
rect 37324 75010 37380 75012
rect 37324 74958 37326 75010
rect 37326 74958 37378 75010
rect 37378 74958 37380 75010
rect 37324 74956 37380 74958
rect 37884 75180 37940 75236
rect 37996 75964 38052 76020
rect 36876 74172 36932 74228
rect 36876 73554 36932 73556
rect 36876 73502 36878 73554
rect 36878 73502 36930 73554
rect 36930 73502 36932 73554
rect 36876 73500 36932 73502
rect 36988 72940 37044 72996
rect 37548 73612 37604 73668
rect 37772 73612 37828 73668
rect 37660 73276 37716 73332
rect 37548 72940 37604 72996
rect 37436 72604 37492 72660
rect 37884 73442 37940 73444
rect 37884 73390 37886 73442
rect 37886 73390 37938 73442
rect 37938 73390 37940 73442
rect 37884 73388 37940 73390
rect 37884 72546 37940 72548
rect 37884 72494 37886 72546
rect 37886 72494 37938 72546
rect 37938 72494 37940 72546
rect 37884 72492 37940 72494
rect 37772 71932 37828 71988
rect 37772 70812 37828 70868
rect 36764 70364 36820 70420
rect 36540 70140 36596 70196
rect 37212 70194 37268 70196
rect 37212 70142 37214 70194
rect 37214 70142 37266 70194
rect 37266 70142 37268 70194
rect 37212 70140 37268 70142
rect 37548 70194 37604 70196
rect 37548 70142 37550 70194
rect 37550 70142 37602 70194
rect 37602 70142 37604 70194
rect 37548 70140 37604 70142
rect 38220 74898 38276 74900
rect 38220 74846 38222 74898
rect 38222 74846 38274 74898
rect 38274 74846 38276 74898
rect 38220 74844 38276 74846
rect 38108 74396 38164 74452
rect 38556 76524 38612 76580
rect 38780 76748 38836 76804
rect 39116 76578 39172 76580
rect 39116 76526 39118 76578
rect 39118 76526 39170 76578
rect 39170 76526 39172 76578
rect 39116 76524 39172 76526
rect 38892 75852 38948 75908
rect 38668 75628 38724 75684
rect 38556 74956 38612 75012
rect 38108 74114 38164 74116
rect 38108 74062 38110 74114
rect 38110 74062 38162 74114
rect 38162 74062 38164 74114
rect 38108 74060 38164 74062
rect 38780 75404 38836 75460
rect 38780 75180 38836 75236
rect 38668 74786 38724 74788
rect 38668 74734 38670 74786
rect 38670 74734 38722 74786
rect 38722 74734 38724 74786
rect 38668 74732 38724 74734
rect 39004 75010 39060 75012
rect 39004 74958 39006 75010
rect 39006 74958 39058 75010
rect 39058 74958 39060 75010
rect 39004 74956 39060 74958
rect 38444 73836 38500 73892
rect 38780 73612 38836 73668
rect 39004 73890 39060 73892
rect 39004 73838 39006 73890
rect 39006 73838 39058 73890
rect 39058 73838 39060 73890
rect 39004 73836 39060 73838
rect 38892 73500 38948 73556
rect 38444 73330 38500 73332
rect 38444 73278 38446 73330
rect 38446 73278 38498 73330
rect 38498 73278 38500 73330
rect 38444 73276 38500 73278
rect 38444 72492 38500 72548
rect 38668 72828 38724 72884
rect 38556 72322 38612 72324
rect 38556 72270 38558 72322
rect 38558 72270 38610 72322
rect 38610 72270 38612 72322
rect 38556 72268 38612 72270
rect 38220 71090 38276 71092
rect 38220 71038 38222 71090
rect 38222 71038 38274 71090
rect 38274 71038 38276 71090
rect 38220 71036 38276 71038
rect 38108 70924 38164 70980
rect 38780 71932 38836 71988
rect 38892 73276 38948 73332
rect 38780 71708 38836 71764
rect 39004 72268 39060 72324
rect 39004 71762 39060 71764
rect 39004 71710 39006 71762
rect 39006 71710 39058 71762
rect 39058 71710 39060 71762
rect 39004 71708 39060 71710
rect 39004 71484 39060 71540
rect 39004 71036 39060 71092
rect 39004 70588 39060 70644
rect 4476 69802 4532 69804
rect 4476 69750 4478 69802
rect 4478 69750 4530 69802
rect 4530 69750 4532 69802
rect 4476 69748 4532 69750
rect 4580 69802 4636 69804
rect 4580 69750 4582 69802
rect 4582 69750 4634 69802
rect 4634 69750 4636 69802
rect 4580 69748 4636 69750
rect 4684 69802 4740 69804
rect 4684 69750 4686 69802
rect 4686 69750 4738 69802
rect 4738 69750 4740 69802
rect 4684 69748 4740 69750
rect 35196 69802 35252 69804
rect 35196 69750 35198 69802
rect 35198 69750 35250 69802
rect 35250 69750 35252 69802
rect 35196 69748 35252 69750
rect 35300 69802 35356 69804
rect 35300 69750 35302 69802
rect 35302 69750 35354 69802
rect 35354 69750 35356 69802
rect 35300 69748 35356 69750
rect 35404 69802 35460 69804
rect 35404 69750 35406 69802
rect 35406 69750 35458 69802
rect 35458 69750 35460 69802
rect 35404 69748 35460 69750
rect 39228 72380 39284 72436
rect 39340 76300 39396 76356
rect 41692 76354 41748 76356
rect 41692 76302 41694 76354
rect 41694 76302 41746 76354
rect 41746 76302 41748 76354
rect 41692 76300 41748 76302
rect 40012 76188 40068 76244
rect 39900 75740 39956 75796
rect 40236 75852 40292 75908
rect 40460 75794 40516 75796
rect 40460 75742 40462 75794
rect 40462 75742 40514 75794
rect 40514 75742 40516 75794
rect 40460 75740 40516 75742
rect 39228 71932 39284 71988
rect 39228 70924 39284 70980
rect 39228 70140 39284 70196
rect 40124 75292 40180 75348
rect 40012 75122 40068 75124
rect 40012 75070 40014 75122
rect 40014 75070 40066 75122
rect 40066 75070 40068 75122
rect 40012 75068 40068 75070
rect 40236 74956 40292 75012
rect 40460 75516 40516 75572
rect 40012 74172 40068 74228
rect 39452 73948 39508 74004
rect 39900 74002 39956 74004
rect 39900 73950 39902 74002
rect 39902 73950 39954 74002
rect 39954 73950 39956 74002
rect 39900 73948 39956 73950
rect 39676 73836 39732 73892
rect 40348 74172 40404 74228
rect 41132 75682 41188 75684
rect 41132 75630 41134 75682
rect 41134 75630 41186 75682
rect 41186 75630 41188 75682
rect 41132 75628 41188 75630
rect 41692 75570 41748 75572
rect 41692 75518 41694 75570
rect 41694 75518 41746 75570
rect 41746 75518 41748 75570
rect 41692 75516 41748 75518
rect 41244 75458 41300 75460
rect 41244 75406 41246 75458
rect 41246 75406 41298 75458
rect 41298 75406 41300 75458
rect 41244 75404 41300 75406
rect 41132 75292 41188 75348
rect 40684 75068 40740 75124
rect 41020 75122 41076 75124
rect 41020 75070 41022 75122
rect 41022 75070 41074 75122
rect 41074 75070 41076 75122
rect 41020 75068 41076 75070
rect 40796 74956 40852 75012
rect 40908 74844 40964 74900
rect 40012 73276 40068 73332
rect 40012 72828 40068 72884
rect 40348 72546 40404 72548
rect 40348 72494 40350 72546
rect 40350 72494 40402 72546
rect 40402 72494 40404 72546
rect 40348 72492 40404 72494
rect 40012 72268 40068 72324
rect 40124 71874 40180 71876
rect 40124 71822 40126 71874
rect 40126 71822 40178 71874
rect 40178 71822 40180 71874
rect 40124 71820 40180 71822
rect 40124 71484 40180 71540
rect 39900 71202 39956 71204
rect 39900 71150 39902 71202
rect 39902 71150 39954 71202
rect 39954 71150 39956 71202
rect 39900 71148 39956 71150
rect 40236 71036 40292 71092
rect 40348 71148 40404 71204
rect 39676 70812 39732 70868
rect 39900 70754 39956 70756
rect 39900 70702 39902 70754
rect 39902 70702 39954 70754
rect 39954 70702 39956 70754
rect 39900 70700 39956 70702
rect 39788 70588 39844 70644
rect 40124 70418 40180 70420
rect 40124 70366 40126 70418
rect 40126 70366 40178 70418
rect 40178 70366 40180 70418
rect 40124 70364 40180 70366
rect 40796 74002 40852 74004
rect 40796 73950 40798 74002
rect 40798 73950 40850 74002
rect 40850 73950 40852 74002
rect 40796 73948 40852 73950
rect 40572 73836 40628 73892
rect 41020 73948 41076 74004
rect 41020 73500 41076 73556
rect 40796 73330 40852 73332
rect 40796 73278 40798 73330
rect 40798 73278 40850 73330
rect 40850 73278 40852 73330
rect 40796 73276 40852 73278
rect 40572 73164 40628 73220
rect 41020 73052 41076 73108
rect 41020 72716 41076 72772
rect 40572 72604 40628 72660
rect 41132 72604 41188 72660
rect 41020 71820 41076 71876
rect 41132 71596 41188 71652
rect 40908 71090 40964 71092
rect 40908 71038 40910 71090
rect 40910 71038 40962 71090
rect 40962 71038 40964 71090
rect 40908 71036 40964 71038
rect 41468 73836 41524 73892
rect 41244 71148 41300 71204
rect 41468 72492 41524 72548
rect 43708 77308 43764 77364
rect 42812 76300 42868 76356
rect 41916 75180 41972 75236
rect 42252 74844 42308 74900
rect 42476 75180 42532 75236
rect 42028 74620 42084 74676
rect 42140 74060 42196 74116
rect 42476 74060 42532 74116
rect 42700 74898 42756 74900
rect 42700 74846 42702 74898
rect 42702 74846 42754 74898
rect 42754 74846 42756 74898
rect 42700 74844 42756 74846
rect 43036 75570 43092 75572
rect 43036 75518 43038 75570
rect 43038 75518 43090 75570
rect 43090 75518 43092 75570
rect 43036 75516 43092 75518
rect 43260 75516 43316 75572
rect 42924 75180 42980 75236
rect 43148 75122 43204 75124
rect 43148 75070 43150 75122
rect 43150 75070 43202 75122
rect 43202 75070 43204 75122
rect 43148 75068 43204 75070
rect 41692 72604 41748 72660
rect 41692 72322 41748 72324
rect 41692 72270 41694 72322
rect 41694 72270 41746 72322
rect 41746 72270 41748 72322
rect 41692 72268 41748 72270
rect 41804 71762 41860 71764
rect 41804 71710 41806 71762
rect 41806 71710 41858 71762
rect 41858 71710 41860 71762
rect 41804 71708 41860 71710
rect 41804 71036 41860 71092
rect 43148 74732 43204 74788
rect 42700 73724 42756 73780
rect 42812 73948 42868 74004
rect 42700 73218 42756 73220
rect 42700 73166 42702 73218
rect 42702 73166 42754 73218
rect 42754 73166 42756 73218
rect 42700 73164 42756 73166
rect 42924 73724 42980 73780
rect 43820 76690 43876 76692
rect 43820 76638 43822 76690
rect 43822 76638 43874 76690
rect 43874 76638 43876 76690
rect 43820 76636 43876 76638
rect 43484 75570 43540 75572
rect 43484 75518 43486 75570
rect 43486 75518 43538 75570
rect 43538 75518 43540 75570
rect 43484 75516 43540 75518
rect 44044 76242 44100 76244
rect 44044 76190 44046 76242
rect 44046 76190 44098 76242
rect 44098 76190 44100 76242
rect 44044 76188 44100 76190
rect 43932 75628 43988 75684
rect 43708 75458 43764 75460
rect 43708 75406 43710 75458
rect 43710 75406 43762 75458
rect 43762 75406 43764 75458
rect 43708 75404 43764 75406
rect 43596 75292 43652 75348
rect 43708 75180 43764 75236
rect 43932 75068 43988 75124
rect 43372 73612 43428 73668
rect 43820 74786 43876 74788
rect 43820 74734 43822 74786
rect 43822 74734 43874 74786
rect 43874 74734 43876 74786
rect 43820 74732 43876 74734
rect 43484 73948 43540 74004
rect 43148 73330 43204 73332
rect 43148 73278 43150 73330
rect 43150 73278 43202 73330
rect 43202 73278 43204 73330
rect 43148 73276 43204 73278
rect 42924 73106 42980 73108
rect 42924 73054 42926 73106
rect 42926 73054 42978 73106
rect 42978 73054 42980 73106
rect 42924 73052 42980 73054
rect 43372 72940 43428 72996
rect 43148 72658 43204 72660
rect 43148 72606 43150 72658
rect 43150 72606 43202 72658
rect 43202 72606 43204 72658
rect 43148 72604 43204 72606
rect 42924 71820 42980 71876
rect 42252 71596 42308 71652
rect 42812 71596 42868 71652
rect 42812 70978 42868 70980
rect 42812 70926 42814 70978
rect 42814 70926 42866 70978
rect 42866 70926 42868 70978
rect 42812 70924 42868 70926
rect 41020 70700 41076 70756
rect 40124 70140 40180 70196
rect 43260 71874 43316 71876
rect 43260 71822 43262 71874
rect 43262 71822 43314 71874
rect 43314 71822 43316 71874
rect 43260 71820 43316 71822
rect 43708 74620 43764 74676
rect 43596 72380 43652 72436
rect 43596 71372 43652 71428
rect 44156 75404 44212 75460
rect 44156 74956 44212 75012
rect 44268 75180 44324 75236
rect 44044 74284 44100 74340
rect 44492 75516 44548 75572
rect 45052 76524 45108 76580
rect 44604 75180 44660 75236
rect 44716 76188 44772 76244
rect 44380 74620 44436 74676
rect 44380 74396 44436 74452
rect 43932 74226 43988 74228
rect 43932 74174 43934 74226
rect 43934 74174 43986 74226
rect 43986 74174 43988 74226
rect 43932 74172 43988 74174
rect 44156 74114 44212 74116
rect 44156 74062 44158 74114
rect 44158 74062 44210 74114
rect 44210 74062 44212 74114
rect 44156 74060 44212 74062
rect 45052 75852 45108 75908
rect 44828 75794 44884 75796
rect 44828 75742 44830 75794
rect 44830 75742 44882 75794
rect 44882 75742 44884 75794
rect 44828 75740 44884 75742
rect 44828 75180 44884 75236
rect 45164 74732 45220 74788
rect 44828 74508 44884 74564
rect 44828 74226 44884 74228
rect 44828 74174 44830 74226
rect 44830 74174 44882 74226
rect 44882 74174 44884 74226
rect 44828 74172 44884 74174
rect 43820 73836 43876 73892
rect 44156 73836 44212 73892
rect 44044 73500 44100 73556
rect 43932 73276 43988 73332
rect 44268 73724 44324 73780
rect 44716 73724 44772 73780
rect 44604 73442 44660 73444
rect 44604 73390 44606 73442
rect 44606 73390 44658 73442
rect 44658 73390 44660 73442
rect 44604 73388 44660 73390
rect 44156 72716 44212 72772
rect 43932 72434 43988 72436
rect 43932 72382 43934 72434
rect 43934 72382 43986 72434
rect 43986 72382 43988 72434
rect 43932 72380 43988 72382
rect 44492 71762 44548 71764
rect 44492 71710 44494 71762
rect 44494 71710 44546 71762
rect 44546 71710 44548 71762
rect 44492 71708 44548 71710
rect 44716 71372 44772 71428
rect 44940 73724 44996 73780
rect 44940 73106 44996 73108
rect 44940 73054 44942 73106
rect 44942 73054 44994 73106
rect 44994 73054 44996 73106
rect 44940 73052 44996 73054
rect 45836 77420 45892 77476
rect 45500 76578 45556 76580
rect 45500 76526 45502 76578
rect 45502 76526 45554 76578
rect 45554 76526 45556 76578
rect 45500 76524 45556 76526
rect 46956 77420 47012 77476
rect 45948 76412 46004 76468
rect 46396 76354 46452 76356
rect 46396 76302 46398 76354
rect 46398 76302 46450 76354
rect 46450 76302 46452 76354
rect 46396 76300 46452 76302
rect 45500 75964 45556 76020
rect 45612 75458 45668 75460
rect 45612 75406 45614 75458
rect 45614 75406 45666 75458
rect 45666 75406 45668 75458
rect 45612 75404 45668 75406
rect 45948 75404 46004 75460
rect 46508 75180 46564 75236
rect 46956 76412 47012 76468
rect 45724 74898 45780 74900
rect 45724 74846 45726 74898
rect 45726 74846 45778 74898
rect 45778 74846 45780 74898
rect 45724 74844 45780 74846
rect 45500 74620 45556 74676
rect 45612 74002 45668 74004
rect 45612 73950 45614 74002
rect 45614 73950 45666 74002
rect 45666 73950 45668 74002
rect 45612 73948 45668 73950
rect 45164 72546 45220 72548
rect 45164 72494 45166 72546
rect 45166 72494 45218 72546
rect 45218 72494 45220 72546
rect 45164 72492 45220 72494
rect 45052 72380 45108 72436
rect 44940 71484 44996 71540
rect 45164 71874 45220 71876
rect 45164 71822 45166 71874
rect 45166 71822 45218 71874
rect 45218 71822 45220 71874
rect 45164 71820 45220 71822
rect 45724 73500 45780 73556
rect 45612 73388 45668 73444
rect 45500 72604 45556 72660
rect 46284 74844 46340 74900
rect 45948 73724 46004 73780
rect 46172 73500 46228 73556
rect 46396 74674 46452 74676
rect 46396 74622 46398 74674
rect 46398 74622 46450 74674
rect 46450 74622 46452 74674
rect 46396 74620 46452 74622
rect 46284 73836 46340 73892
rect 46060 73276 46116 73332
rect 45052 71036 45108 71092
rect 44828 70924 44884 70980
rect 46284 73276 46340 73332
rect 46284 73052 46340 73108
rect 46396 72434 46452 72436
rect 46396 72382 46398 72434
rect 46398 72382 46450 72434
rect 46450 72382 46452 72434
rect 46396 72380 46452 72382
rect 46284 72268 46340 72324
rect 45612 71090 45668 71092
rect 45612 71038 45614 71090
rect 45614 71038 45666 71090
rect 45666 71038 45668 71090
rect 45612 71036 45668 71038
rect 45276 70476 45332 70532
rect 46060 71148 46116 71204
rect 46620 73612 46676 73668
rect 46620 72546 46676 72548
rect 46620 72494 46622 72546
rect 46622 72494 46674 72546
rect 46674 72494 46676 72546
rect 46620 72492 46676 72494
rect 46844 73052 46900 73108
rect 47180 75404 47236 75460
rect 47404 75570 47460 75572
rect 47404 75518 47406 75570
rect 47406 75518 47458 75570
rect 47458 75518 47460 75570
rect 47404 75516 47460 75518
rect 47292 74060 47348 74116
rect 47404 75292 47460 75348
rect 47068 73948 47124 74004
rect 47180 73442 47236 73444
rect 47180 73390 47182 73442
rect 47182 73390 47234 73442
rect 47234 73390 47236 73442
rect 47180 73388 47236 73390
rect 47068 73276 47124 73332
rect 47180 73164 47236 73220
rect 46508 71932 46564 71988
rect 47292 72492 47348 72548
rect 46396 71148 46452 71204
rect 46172 70924 46228 70980
rect 46172 70418 46228 70420
rect 46172 70366 46174 70418
rect 46174 70366 46226 70418
rect 46226 70366 46228 70418
rect 46172 70364 46228 70366
rect 47852 74226 47908 74228
rect 47852 74174 47854 74226
rect 47854 74174 47906 74226
rect 47906 74174 47908 74226
rect 47852 74172 47908 74174
rect 47852 73948 47908 74004
rect 48524 76524 48580 76580
rect 48412 75964 48468 76020
rect 48300 75458 48356 75460
rect 48300 75406 48302 75458
rect 48302 75406 48354 75458
rect 48354 75406 48356 75458
rect 48300 75404 48356 75406
rect 47852 73554 47908 73556
rect 47852 73502 47854 73554
rect 47854 73502 47906 73554
rect 47906 73502 47908 73554
rect 47852 73500 47908 73502
rect 47628 72322 47684 72324
rect 47628 72270 47630 72322
rect 47630 72270 47682 72322
rect 47682 72270 47684 72322
rect 47628 72268 47684 72270
rect 47740 72492 47796 72548
rect 47852 71932 47908 71988
rect 49084 76300 49140 76356
rect 48972 76076 49028 76132
rect 49084 75740 49140 75796
rect 49084 75404 49140 75460
rect 48636 74956 48692 75012
rect 48748 75068 48804 75124
rect 48524 74060 48580 74116
rect 48636 73890 48692 73892
rect 48636 73838 48638 73890
rect 48638 73838 48690 73890
rect 48690 73838 48692 73890
rect 48636 73836 48692 73838
rect 48860 73388 48916 73444
rect 48412 72492 48468 72548
rect 48076 71986 48132 71988
rect 48076 71934 48078 71986
rect 48078 71934 48130 71986
rect 48130 71934 48132 71986
rect 48076 71932 48132 71934
rect 50652 76972 50708 77028
rect 50556 76858 50612 76860
rect 50556 76806 50558 76858
rect 50558 76806 50610 76858
rect 50610 76806 50612 76858
rect 50556 76804 50612 76806
rect 50660 76858 50716 76860
rect 50660 76806 50662 76858
rect 50662 76806 50714 76858
rect 50714 76806 50716 76858
rect 50660 76804 50716 76806
rect 50764 76858 50820 76860
rect 50764 76806 50766 76858
rect 50766 76806 50818 76858
rect 50818 76806 50820 76858
rect 50764 76804 50820 76806
rect 49756 75458 49812 75460
rect 49756 75406 49758 75458
rect 49758 75406 49810 75458
rect 49810 75406 49812 75458
rect 49756 75404 49812 75406
rect 49308 74338 49364 74340
rect 49308 74286 49310 74338
rect 49310 74286 49362 74338
rect 49362 74286 49364 74338
rect 49308 74284 49364 74286
rect 49420 73388 49476 73444
rect 49532 74956 49588 75012
rect 49420 73218 49476 73220
rect 49420 73166 49422 73218
rect 49422 73166 49474 73218
rect 49474 73166 49476 73218
rect 49420 73164 49476 73166
rect 48412 71260 48468 71316
rect 47852 71090 47908 71092
rect 47852 71038 47854 71090
rect 47854 71038 47906 71090
rect 47906 71038 47908 71090
rect 47852 71036 47908 71038
rect 48748 71090 48804 71092
rect 48748 71038 48750 71090
rect 48750 71038 48802 71090
rect 48802 71038 48804 71090
rect 48748 71036 48804 71038
rect 49308 71090 49364 71092
rect 49308 71038 49310 71090
rect 49310 71038 49362 71090
rect 49362 71038 49364 71090
rect 49308 71036 49364 71038
rect 48300 70364 48356 70420
rect 49644 73276 49700 73332
rect 49756 74060 49812 74116
rect 49644 72604 49700 72660
rect 49868 74002 49924 74004
rect 49868 73950 49870 74002
rect 49870 73950 49922 74002
rect 49922 73950 49924 74002
rect 49868 73948 49924 73950
rect 50092 74172 50148 74228
rect 49980 73836 50036 73892
rect 49868 72828 49924 72884
rect 50092 72492 50148 72548
rect 49868 72268 49924 72324
rect 50316 75068 50372 75124
rect 50316 74898 50372 74900
rect 50316 74846 50318 74898
rect 50318 74846 50370 74898
rect 50370 74846 50372 74898
rect 50316 74844 50372 74846
rect 50316 73948 50372 74004
rect 50556 75290 50612 75292
rect 50556 75238 50558 75290
rect 50558 75238 50610 75290
rect 50610 75238 50612 75290
rect 50556 75236 50612 75238
rect 50660 75290 50716 75292
rect 50660 75238 50662 75290
rect 50662 75238 50714 75290
rect 50714 75238 50716 75290
rect 50660 75236 50716 75238
rect 50764 75290 50820 75292
rect 50764 75238 50766 75290
rect 50766 75238 50818 75290
rect 50818 75238 50820 75290
rect 50764 75236 50820 75238
rect 50764 74956 50820 75012
rect 50988 75068 51044 75124
rect 50876 74844 50932 74900
rect 50652 74114 50708 74116
rect 50652 74062 50654 74114
rect 50654 74062 50706 74114
rect 50706 74062 50708 74114
rect 50652 74060 50708 74062
rect 50876 74002 50932 74004
rect 50876 73950 50878 74002
rect 50878 73950 50930 74002
rect 50930 73950 50932 74002
rect 50876 73948 50932 73950
rect 50556 73722 50612 73724
rect 50556 73670 50558 73722
rect 50558 73670 50610 73722
rect 50610 73670 50612 73722
rect 50556 73668 50612 73670
rect 50660 73722 50716 73724
rect 50660 73670 50662 73722
rect 50662 73670 50714 73722
rect 50714 73670 50716 73722
rect 50660 73668 50716 73670
rect 50764 73722 50820 73724
rect 50764 73670 50766 73722
rect 50766 73670 50818 73722
rect 50818 73670 50820 73722
rect 50764 73668 50820 73670
rect 51100 74284 51156 74340
rect 51548 76972 51604 77028
rect 51436 74898 51492 74900
rect 51436 74846 51438 74898
rect 51438 74846 51490 74898
rect 51490 74846 51492 74898
rect 51436 74844 51492 74846
rect 51996 76412 52052 76468
rect 53228 77196 53284 77252
rect 52892 76972 52948 77028
rect 52668 76300 52724 76356
rect 52332 75964 52388 76020
rect 53116 75906 53172 75908
rect 53116 75854 53118 75906
rect 53118 75854 53170 75906
rect 53170 75854 53172 75906
rect 53116 75852 53172 75854
rect 53004 75682 53060 75684
rect 53004 75630 53006 75682
rect 53006 75630 53058 75682
rect 53058 75630 53060 75682
rect 53004 75628 53060 75630
rect 51660 75180 51716 75236
rect 51548 74732 51604 74788
rect 51212 74060 51268 74116
rect 51324 74172 51380 74228
rect 51436 74060 51492 74116
rect 51100 74002 51156 74004
rect 51100 73950 51102 74002
rect 51102 73950 51154 74002
rect 51154 73950 51156 74002
rect 51100 73948 51156 73950
rect 51548 73612 51604 73668
rect 51996 74844 52052 74900
rect 51884 74060 51940 74116
rect 51996 74508 52052 74564
rect 52108 74284 52164 74340
rect 53004 75010 53060 75012
rect 53004 74958 53006 75010
rect 53006 74958 53058 75010
rect 53058 74958 53060 75010
rect 53004 74956 53060 74958
rect 52892 74620 52948 74676
rect 52780 74172 52836 74228
rect 51772 73890 51828 73892
rect 51772 73838 51774 73890
rect 51774 73838 51826 73890
rect 51826 73838 51828 73890
rect 51772 73836 51828 73838
rect 50316 73276 50372 73332
rect 50764 73218 50820 73220
rect 50764 73166 50766 73218
rect 50766 73166 50818 73218
rect 50818 73166 50820 73218
rect 50764 73164 50820 73166
rect 50876 72716 50932 72772
rect 50764 72546 50820 72548
rect 50764 72494 50766 72546
rect 50766 72494 50818 72546
rect 50818 72494 50820 72546
rect 50764 72492 50820 72494
rect 50316 72268 50372 72324
rect 50988 72268 51044 72324
rect 51100 73052 51156 73108
rect 50556 72154 50612 72156
rect 50556 72102 50558 72154
rect 50558 72102 50610 72154
rect 50610 72102 50612 72154
rect 50556 72100 50612 72102
rect 50660 72154 50716 72156
rect 50660 72102 50662 72154
rect 50662 72102 50714 72154
rect 50714 72102 50716 72154
rect 50660 72100 50716 72102
rect 50764 72154 50820 72156
rect 50764 72102 50766 72154
rect 50766 72102 50818 72154
rect 50818 72102 50820 72154
rect 50764 72100 50820 72102
rect 50204 71762 50260 71764
rect 50204 71710 50206 71762
rect 50206 71710 50258 71762
rect 50258 71710 50260 71762
rect 50204 71708 50260 71710
rect 51548 72658 51604 72660
rect 51548 72606 51550 72658
rect 51550 72606 51602 72658
rect 51602 72606 51604 72658
rect 51548 72604 51604 72606
rect 54012 77308 54068 77364
rect 53340 76636 53396 76692
rect 53900 76578 53956 76580
rect 53900 76526 53902 76578
rect 53902 76526 53954 76578
rect 53954 76526 53956 76578
rect 53900 76524 53956 76526
rect 54236 76300 54292 76356
rect 54348 75964 54404 76020
rect 53564 75740 53620 75796
rect 54124 75682 54180 75684
rect 54124 75630 54126 75682
rect 54126 75630 54178 75682
rect 54178 75630 54180 75682
rect 54124 75628 54180 75630
rect 53788 75570 53844 75572
rect 53788 75518 53790 75570
rect 53790 75518 53842 75570
rect 53842 75518 53844 75570
rect 53788 75516 53844 75518
rect 51996 73388 52052 73444
rect 52332 73612 52388 73668
rect 51772 72716 51828 72772
rect 51996 72604 52052 72660
rect 51884 72546 51940 72548
rect 51884 72494 51886 72546
rect 51886 72494 51938 72546
rect 51938 72494 51940 72546
rect 51884 72492 51940 72494
rect 50876 71090 50932 71092
rect 50876 71038 50878 71090
rect 50878 71038 50930 71090
rect 50930 71038 50932 71090
rect 50876 71036 50932 71038
rect 51548 72268 51604 72324
rect 50556 70586 50612 70588
rect 50556 70534 50558 70586
rect 50558 70534 50610 70586
rect 50610 70534 50612 70586
rect 50556 70532 50612 70534
rect 50660 70586 50716 70588
rect 50660 70534 50662 70586
rect 50662 70534 50714 70586
rect 50714 70534 50716 70586
rect 50660 70532 50716 70534
rect 50764 70586 50820 70588
rect 50764 70534 50766 70586
rect 50766 70534 50818 70586
rect 50818 70534 50820 70586
rect 50764 70532 50820 70534
rect 50204 70418 50260 70420
rect 50204 70366 50206 70418
rect 50206 70366 50258 70418
rect 50258 70366 50260 70418
rect 50204 70364 50260 70366
rect 50652 70418 50708 70420
rect 50652 70366 50654 70418
rect 50654 70366 50706 70418
rect 50706 70366 50708 70418
rect 50652 70364 50708 70366
rect 52108 72492 52164 72548
rect 51884 71708 51940 71764
rect 53116 73388 53172 73444
rect 52444 72546 52500 72548
rect 52444 72494 52446 72546
rect 52446 72494 52498 72546
rect 52498 72494 52500 72546
rect 52444 72492 52500 72494
rect 53004 72492 53060 72548
rect 52668 72434 52724 72436
rect 52668 72382 52670 72434
rect 52670 72382 52722 72434
rect 52722 72382 52724 72434
rect 52668 72380 52724 72382
rect 52892 72268 52948 72324
rect 53788 74284 53844 74340
rect 54012 75458 54068 75460
rect 54012 75406 54014 75458
rect 54014 75406 54066 75458
rect 54066 75406 54068 75458
rect 54012 75404 54068 75406
rect 54460 75682 54516 75684
rect 54460 75630 54462 75682
rect 54462 75630 54514 75682
rect 54514 75630 54516 75682
rect 54460 75628 54516 75630
rect 54012 74956 54068 75012
rect 53676 74172 53732 74228
rect 54348 74898 54404 74900
rect 54348 74846 54350 74898
rect 54350 74846 54402 74898
rect 54402 74846 54404 74898
rect 54348 74844 54404 74846
rect 54124 73500 54180 73556
rect 53564 72716 53620 72772
rect 53340 72604 53396 72660
rect 53228 72492 53284 72548
rect 54124 72268 54180 72324
rect 52556 70476 52612 70532
rect 51660 70418 51716 70420
rect 51660 70366 51662 70418
rect 51662 70366 51714 70418
rect 51714 70366 51716 70418
rect 51660 70364 51716 70366
rect 54796 75180 54852 75236
rect 55132 75682 55188 75684
rect 55132 75630 55134 75682
rect 55134 75630 55186 75682
rect 55186 75630 55188 75682
rect 55132 75628 55188 75630
rect 55020 75458 55076 75460
rect 55020 75406 55022 75458
rect 55022 75406 55074 75458
rect 55074 75406 55076 75458
rect 55020 75404 55076 75406
rect 55020 75180 55076 75236
rect 54460 73836 54516 73892
rect 54572 74284 54628 74340
rect 54684 74114 54740 74116
rect 54684 74062 54686 74114
rect 54686 74062 54738 74114
rect 54738 74062 54740 74114
rect 54684 74060 54740 74062
rect 54460 72716 54516 72772
rect 54348 72434 54404 72436
rect 54348 72382 54350 72434
rect 54350 72382 54402 72434
rect 54402 72382 54404 72434
rect 54348 72380 54404 72382
rect 53004 70418 53060 70420
rect 53004 70366 53006 70418
rect 53006 70366 53058 70418
rect 53058 70366 53060 70418
rect 53004 70364 53060 70366
rect 54684 72546 54740 72548
rect 54684 72494 54686 72546
rect 54686 72494 54738 72546
rect 54738 72494 54740 72546
rect 54684 72492 54740 72494
rect 54572 70476 54628 70532
rect 54236 70418 54292 70420
rect 54236 70366 54238 70418
rect 54238 70366 54290 70418
rect 54290 70366 54292 70418
rect 54236 70364 54292 70366
rect 54124 70252 54180 70308
rect 53452 70082 53508 70084
rect 53452 70030 53454 70082
rect 53454 70030 53506 70082
rect 53506 70030 53508 70082
rect 53452 70028 53508 70030
rect 55244 75180 55300 75236
rect 55356 75068 55412 75124
rect 55580 75516 55636 75572
rect 54908 73890 54964 73892
rect 54908 73838 54910 73890
rect 54910 73838 54962 73890
rect 54962 73838 54964 73890
rect 54908 73836 54964 73838
rect 54908 73442 54964 73444
rect 54908 73390 54910 73442
rect 54910 73390 54962 73442
rect 54962 73390 54964 73442
rect 54908 73388 54964 73390
rect 54908 72716 54964 72772
rect 55468 74674 55524 74676
rect 55468 74622 55470 74674
rect 55470 74622 55522 74674
rect 55522 74622 55524 74674
rect 55468 74620 55524 74622
rect 55356 73836 55412 73892
rect 55356 73554 55412 73556
rect 55356 73502 55358 73554
rect 55358 73502 55410 73554
rect 55410 73502 55412 73554
rect 55356 73500 55412 73502
rect 56588 77532 56644 77588
rect 56140 75852 56196 75908
rect 56140 75458 56196 75460
rect 56140 75406 56142 75458
rect 56142 75406 56194 75458
rect 56194 75406 56196 75458
rect 56140 75404 56196 75406
rect 56028 75292 56084 75348
rect 55804 75180 55860 75236
rect 55692 74844 55748 74900
rect 55692 74284 55748 74340
rect 55692 73164 55748 73220
rect 56028 74002 56084 74004
rect 56028 73950 56030 74002
rect 56030 73950 56082 74002
rect 56082 73950 56084 74002
rect 56028 73948 56084 73950
rect 56028 73554 56084 73556
rect 56028 73502 56030 73554
rect 56030 73502 56082 73554
rect 56082 73502 56084 73554
rect 56028 73500 56084 73502
rect 55916 73388 55972 73444
rect 56364 75852 56420 75908
rect 56476 75570 56532 75572
rect 56476 75518 56478 75570
rect 56478 75518 56530 75570
rect 56530 75518 56532 75570
rect 56476 75516 56532 75518
rect 56700 76524 56756 76580
rect 57932 76578 57988 76580
rect 57932 76526 57934 76578
rect 57934 76526 57986 76578
rect 57986 76526 57988 76578
rect 57932 76524 57988 76526
rect 56924 75852 56980 75908
rect 57036 75180 57092 75236
rect 56588 74172 56644 74228
rect 56924 74060 56980 74116
rect 57036 74620 57092 74676
rect 56252 73164 56308 73220
rect 55244 71820 55300 71876
rect 55468 70924 55524 70980
rect 55244 70700 55300 70756
rect 55468 70754 55524 70756
rect 55468 70702 55470 70754
rect 55470 70702 55522 70754
rect 55522 70702 55524 70754
rect 55468 70700 55524 70702
rect 55356 70476 55412 70532
rect 56588 73052 56644 73108
rect 56140 71202 56196 71204
rect 56140 71150 56142 71202
rect 56142 71150 56194 71202
rect 56194 71150 56196 71202
rect 56140 71148 56196 71150
rect 57372 75180 57428 75236
rect 57148 73836 57204 73892
rect 60620 77308 60676 77364
rect 58604 76524 58660 76580
rect 58380 76076 58436 76132
rect 58044 75404 58100 75460
rect 57596 74114 57652 74116
rect 57596 74062 57598 74114
rect 57598 74062 57650 74114
rect 57650 74062 57652 74114
rect 57596 74060 57652 74062
rect 58044 75180 58100 75236
rect 57932 74002 57988 74004
rect 57932 73950 57934 74002
rect 57934 73950 57986 74002
rect 57986 73950 57988 74002
rect 57932 73948 57988 73950
rect 57484 73724 57540 73780
rect 56924 73276 56980 73332
rect 56812 73164 56868 73220
rect 57148 72604 57204 72660
rect 57820 73500 57876 73556
rect 58268 74956 58324 75012
rect 58268 74508 58324 74564
rect 58940 75740 58996 75796
rect 59164 75852 59220 75908
rect 58940 75068 58996 75124
rect 59836 76412 59892 76468
rect 59612 75964 59668 76020
rect 59948 75570 60004 75572
rect 59948 75518 59950 75570
rect 59950 75518 60002 75570
rect 60002 75518 60004 75570
rect 59948 75516 60004 75518
rect 58828 74956 58884 75012
rect 58828 74732 58884 74788
rect 59164 74898 59220 74900
rect 59164 74846 59166 74898
rect 59166 74846 59218 74898
rect 59218 74846 59220 74898
rect 59164 74844 59220 74846
rect 59164 74172 59220 74228
rect 58604 73724 58660 73780
rect 57708 73330 57764 73332
rect 57708 73278 57710 73330
rect 57710 73278 57762 73330
rect 57762 73278 57764 73330
rect 57708 73276 57764 73278
rect 57484 72604 57540 72660
rect 57036 72380 57092 72436
rect 55916 70978 55972 70980
rect 55916 70926 55918 70978
rect 55918 70926 55970 70978
rect 55970 70926 55972 70978
rect 55916 70924 55972 70926
rect 55580 70364 55636 70420
rect 56028 70418 56084 70420
rect 56028 70366 56030 70418
rect 56030 70366 56082 70418
rect 56082 70366 56084 70418
rect 56028 70364 56084 70366
rect 56476 70418 56532 70420
rect 56476 70366 56478 70418
rect 56478 70366 56530 70418
rect 56530 70366 56532 70418
rect 56476 70364 56532 70366
rect 56700 72044 56756 72100
rect 56700 71874 56756 71876
rect 56700 71822 56702 71874
rect 56702 71822 56754 71874
rect 56754 71822 56756 71874
rect 56700 71820 56756 71822
rect 57372 71820 57428 71876
rect 57932 71874 57988 71876
rect 57932 71822 57934 71874
rect 57934 71822 57986 71874
rect 57986 71822 57988 71874
rect 57932 71820 57988 71822
rect 57372 71202 57428 71204
rect 57372 71150 57374 71202
rect 57374 71150 57426 71202
rect 57426 71150 57428 71202
rect 57372 71148 57428 71150
rect 58828 72492 58884 72548
rect 58716 72044 58772 72100
rect 59276 73330 59332 73332
rect 59276 73278 59278 73330
rect 59278 73278 59330 73330
rect 59330 73278 59332 73330
rect 59276 73276 59332 73278
rect 59500 74284 59556 74340
rect 59836 75180 59892 75236
rect 59724 74956 59780 75012
rect 59948 74956 60004 75012
rect 59724 74508 59780 74564
rect 60508 76690 60564 76692
rect 60508 76638 60510 76690
rect 60510 76638 60562 76690
rect 60562 76638 60564 76690
rect 60508 76636 60564 76638
rect 61628 75628 61684 75684
rect 61404 75516 61460 75572
rect 61740 75292 61796 75348
rect 60172 75180 60228 75236
rect 61628 75068 61684 75124
rect 60172 75010 60228 75012
rect 60172 74958 60174 75010
rect 60174 74958 60226 75010
rect 60226 74958 60228 75010
rect 60172 74956 60228 74958
rect 61852 74956 61908 75012
rect 61516 74898 61572 74900
rect 61516 74846 61518 74898
rect 61518 74846 61570 74898
rect 61570 74846 61572 74898
rect 61516 74844 61572 74846
rect 60284 74786 60340 74788
rect 60284 74734 60286 74786
rect 60286 74734 60338 74786
rect 60338 74734 60340 74786
rect 60284 74732 60340 74734
rect 60844 74674 60900 74676
rect 60844 74622 60846 74674
rect 60846 74622 60898 74674
rect 60898 74622 60900 74674
rect 60844 74620 60900 74622
rect 60956 74508 61012 74564
rect 61404 74732 61460 74788
rect 60620 74284 60676 74340
rect 60508 73890 60564 73892
rect 60508 73838 60510 73890
rect 60510 73838 60562 73890
rect 60562 73838 60564 73890
rect 60508 73836 60564 73838
rect 59836 73612 59892 73668
rect 59276 73052 59332 73108
rect 60172 73276 60228 73332
rect 59164 72434 59220 72436
rect 59164 72382 59166 72434
rect 59166 72382 59218 72434
rect 59218 72382 59220 72434
rect 59164 72380 59220 72382
rect 59276 71986 59332 71988
rect 59276 71934 59278 71986
rect 59278 71934 59330 71986
rect 59330 71934 59332 71986
rect 59276 71932 59332 71934
rect 59724 72658 59780 72660
rect 59724 72606 59726 72658
rect 59726 72606 59778 72658
rect 59778 72606 59780 72658
rect 59724 72604 59780 72606
rect 61628 74284 61684 74340
rect 61404 74060 61460 74116
rect 60956 73724 61012 73780
rect 60396 72044 60452 72100
rect 62748 76524 62804 76580
rect 63532 76524 63588 76580
rect 62412 76466 62468 76468
rect 62412 76414 62414 76466
rect 62414 76414 62466 76466
rect 62466 76414 62468 76466
rect 62412 76412 62468 76414
rect 62860 76242 62916 76244
rect 62860 76190 62862 76242
rect 62862 76190 62914 76242
rect 62914 76190 62916 76242
rect 62860 76188 62916 76190
rect 62524 76076 62580 76132
rect 62412 75458 62468 75460
rect 62412 75406 62414 75458
rect 62414 75406 62466 75458
rect 62466 75406 62468 75458
rect 62412 75404 62468 75406
rect 62076 75068 62132 75124
rect 62188 75180 62244 75236
rect 63084 75570 63140 75572
rect 63084 75518 63086 75570
rect 63086 75518 63138 75570
rect 63138 75518 63140 75570
rect 63084 75516 63140 75518
rect 62860 75122 62916 75124
rect 62860 75070 62862 75122
rect 62862 75070 62914 75122
rect 62914 75070 62916 75122
rect 62860 75068 62916 75070
rect 63420 74786 63476 74788
rect 63420 74734 63422 74786
rect 63422 74734 63474 74786
rect 63474 74734 63476 74786
rect 63420 74732 63476 74734
rect 61964 74172 62020 74228
rect 62972 74226 63028 74228
rect 62972 74174 62974 74226
rect 62974 74174 63026 74226
rect 63026 74174 63028 74226
rect 62972 74172 63028 74174
rect 63868 75516 63924 75572
rect 64988 76578 65044 76580
rect 64988 76526 64990 76578
rect 64990 76526 65042 76578
rect 65042 76526 65044 76578
rect 64988 76524 65044 76526
rect 65212 76524 65268 76580
rect 63868 74956 63924 75012
rect 65916 76074 65972 76076
rect 65916 76022 65918 76074
rect 65918 76022 65970 76074
rect 65970 76022 65972 76074
rect 65916 76020 65972 76022
rect 66020 76074 66076 76076
rect 66020 76022 66022 76074
rect 66022 76022 66074 76074
rect 66074 76022 66076 76074
rect 66020 76020 66076 76022
rect 66124 76074 66180 76076
rect 66124 76022 66126 76074
rect 66126 76022 66178 76074
rect 66178 76022 66180 76074
rect 66124 76020 66180 76022
rect 66780 75516 66836 75572
rect 65916 74506 65972 74508
rect 65916 74454 65918 74506
rect 65918 74454 65970 74506
rect 65970 74454 65972 74506
rect 65916 74452 65972 74454
rect 66020 74506 66076 74508
rect 66020 74454 66022 74506
rect 66022 74454 66074 74506
rect 66074 74454 66076 74506
rect 66020 74452 66076 74454
rect 66124 74506 66180 74508
rect 66124 74454 66126 74506
rect 66126 74454 66178 74506
rect 66178 74454 66180 74506
rect 66124 74452 66180 74454
rect 65772 74284 65828 74340
rect 62076 74114 62132 74116
rect 62076 74062 62078 74114
rect 62078 74062 62130 74114
rect 62130 74062 62132 74114
rect 62076 74060 62132 74062
rect 68796 76748 68852 76804
rect 69356 76748 69412 76804
rect 68124 76636 68180 76692
rect 68012 76578 68068 76580
rect 68012 76526 68014 76578
rect 68014 76526 68066 76578
rect 68066 76526 68068 76578
rect 68012 76524 68068 76526
rect 69020 76300 69076 76356
rect 69020 75570 69076 75572
rect 69020 75518 69022 75570
rect 69022 75518 69074 75570
rect 69074 75518 69076 75570
rect 69020 75516 69076 75518
rect 69916 76690 69972 76692
rect 69916 76638 69918 76690
rect 69918 76638 69970 76690
rect 69970 76638 69972 76690
rect 69916 76636 69972 76638
rect 70476 76748 70532 76804
rect 70924 77420 70980 77476
rect 70812 76524 70868 76580
rect 70140 75516 70196 75572
rect 70700 75570 70756 75572
rect 70700 75518 70702 75570
rect 70702 75518 70754 75570
rect 70754 75518 70756 75570
rect 70700 75516 70756 75518
rect 69468 75404 69524 75460
rect 70028 75458 70084 75460
rect 70028 75406 70030 75458
rect 70030 75406 70082 75458
rect 70082 75406 70084 75458
rect 70028 75404 70084 75406
rect 73052 76578 73108 76580
rect 73052 76526 73054 76578
rect 73054 76526 73106 76578
rect 73106 76526 73108 76578
rect 73052 76524 73108 76526
rect 72828 75404 72884 75460
rect 66892 73276 66948 73332
rect 65916 72938 65972 72940
rect 65916 72886 65918 72938
rect 65918 72886 65970 72938
rect 65970 72886 65972 72938
rect 65916 72884 65972 72886
rect 66020 72938 66076 72940
rect 66020 72886 66022 72938
rect 66022 72886 66074 72938
rect 66074 72886 66076 72938
rect 66020 72884 66076 72886
rect 66124 72938 66180 72940
rect 66124 72886 66126 72938
rect 66126 72886 66178 72938
rect 66178 72886 66180 72938
rect 66124 72884 66180 72886
rect 61404 71932 61460 71988
rect 58940 71820 58996 71876
rect 65916 71370 65972 71372
rect 65916 71318 65918 71370
rect 65918 71318 65970 71370
rect 65970 71318 65972 71370
rect 65916 71316 65972 71318
rect 66020 71370 66076 71372
rect 66020 71318 66022 71370
rect 66022 71318 66074 71370
rect 66074 71318 66076 71370
rect 66020 71316 66076 71318
rect 66124 71370 66180 71372
rect 66124 71318 66126 71370
rect 66126 71318 66178 71370
rect 66178 71318 66180 71370
rect 66124 71316 66180 71318
rect 73500 75516 73556 75572
rect 73948 75570 74004 75572
rect 73948 75518 73950 75570
rect 73950 75518 74002 75570
rect 74002 75518 74004 75570
rect 73948 75516 74004 75518
rect 73388 75404 73444 75460
rect 74508 76242 74564 76244
rect 74508 76190 74510 76242
rect 74510 76190 74562 76242
rect 74562 76190 74564 76242
rect 74508 76188 74564 76190
rect 75068 75628 75124 75684
rect 74956 75516 75012 75572
rect 76972 75570 77028 75572
rect 76972 75518 76974 75570
rect 76974 75518 77026 75570
rect 77026 75518 77028 75570
rect 76972 75516 77028 75518
rect 77420 75516 77476 75572
rect 77644 74172 77700 74228
rect 78092 74226 78148 74228
rect 78092 74174 78094 74226
rect 78094 74174 78146 74226
rect 78146 74174 78148 74226
rect 78092 74172 78148 74174
rect 73052 71036 73108 71092
rect 57036 70978 57092 70980
rect 57036 70926 57038 70978
rect 57038 70926 57090 70978
rect 57090 70926 57092 70978
rect 57036 70924 57092 70926
rect 56588 70252 56644 70308
rect 56924 70306 56980 70308
rect 56924 70254 56926 70306
rect 56926 70254 56978 70306
rect 56978 70254 56980 70306
rect 56924 70252 56980 70254
rect 55580 70028 55636 70084
rect 65916 69802 65972 69804
rect 65916 69750 65918 69802
rect 65918 69750 65970 69802
rect 65970 69750 65972 69802
rect 65916 69748 65972 69750
rect 66020 69802 66076 69804
rect 66020 69750 66022 69802
rect 66022 69750 66074 69802
rect 66074 69750 66076 69802
rect 66020 69748 66076 69750
rect 66124 69802 66180 69804
rect 66124 69750 66126 69802
rect 66126 69750 66178 69802
rect 66178 69750 66180 69802
rect 66124 69748 66180 69750
rect 19836 69018 19892 69020
rect 19836 68966 19838 69018
rect 19838 68966 19890 69018
rect 19890 68966 19892 69018
rect 19836 68964 19892 68966
rect 19940 69018 19996 69020
rect 19940 68966 19942 69018
rect 19942 68966 19994 69018
rect 19994 68966 19996 69018
rect 19940 68964 19996 68966
rect 20044 69018 20100 69020
rect 20044 68966 20046 69018
rect 20046 68966 20098 69018
rect 20098 68966 20100 69018
rect 20044 68964 20100 68966
rect 50556 69018 50612 69020
rect 50556 68966 50558 69018
rect 50558 68966 50610 69018
rect 50610 68966 50612 69018
rect 50556 68964 50612 68966
rect 50660 69018 50716 69020
rect 50660 68966 50662 69018
rect 50662 68966 50714 69018
rect 50714 68966 50716 69018
rect 50660 68964 50716 68966
rect 50764 69018 50820 69020
rect 50764 68966 50766 69018
rect 50766 68966 50818 69018
rect 50818 68966 50820 69018
rect 50764 68964 50820 68966
rect 4476 68234 4532 68236
rect 4476 68182 4478 68234
rect 4478 68182 4530 68234
rect 4530 68182 4532 68234
rect 4476 68180 4532 68182
rect 4580 68234 4636 68236
rect 4580 68182 4582 68234
rect 4582 68182 4634 68234
rect 4634 68182 4636 68234
rect 4580 68180 4636 68182
rect 4684 68234 4740 68236
rect 4684 68182 4686 68234
rect 4686 68182 4738 68234
rect 4738 68182 4740 68234
rect 4684 68180 4740 68182
rect 35196 68234 35252 68236
rect 35196 68182 35198 68234
rect 35198 68182 35250 68234
rect 35250 68182 35252 68234
rect 35196 68180 35252 68182
rect 35300 68234 35356 68236
rect 35300 68182 35302 68234
rect 35302 68182 35354 68234
rect 35354 68182 35356 68234
rect 35300 68180 35356 68182
rect 35404 68234 35460 68236
rect 35404 68182 35406 68234
rect 35406 68182 35458 68234
rect 35458 68182 35460 68234
rect 35404 68180 35460 68182
rect 65916 68234 65972 68236
rect 65916 68182 65918 68234
rect 65918 68182 65970 68234
rect 65970 68182 65972 68234
rect 65916 68180 65972 68182
rect 66020 68234 66076 68236
rect 66020 68182 66022 68234
rect 66022 68182 66074 68234
rect 66074 68182 66076 68234
rect 66020 68180 66076 68182
rect 66124 68234 66180 68236
rect 66124 68182 66126 68234
rect 66126 68182 66178 68234
rect 66178 68182 66180 68234
rect 66124 68180 66180 68182
rect 19836 67450 19892 67452
rect 19836 67398 19838 67450
rect 19838 67398 19890 67450
rect 19890 67398 19892 67450
rect 19836 67396 19892 67398
rect 19940 67450 19996 67452
rect 19940 67398 19942 67450
rect 19942 67398 19994 67450
rect 19994 67398 19996 67450
rect 19940 67396 19996 67398
rect 20044 67450 20100 67452
rect 20044 67398 20046 67450
rect 20046 67398 20098 67450
rect 20098 67398 20100 67450
rect 20044 67396 20100 67398
rect 50556 67450 50612 67452
rect 50556 67398 50558 67450
rect 50558 67398 50610 67450
rect 50610 67398 50612 67450
rect 50556 67396 50612 67398
rect 50660 67450 50716 67452
rect 50660 67398 50662 67450
rect 50662 67398 50714 67450
rect 50714 67398 50716 67450
rect 50660 67396 50716 67398
rect 50764 67450 50820 67452
rect 50764 67398 50766 67450
rect 50766 67398 50818 67450
rect 50818 67398 50820 67450
rect 50764 67396 50820 67398
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 35196 66666 35252 66668
rect 35196 66614 35198 66666
rect 35198 66614 35250 66666
rect 35250 66614 35252 66666
rect 35196 66612 35252 66614
rect 35300 66666 35356 66668
rect 35300 66614 35302 66666
rect 35302 66614 35354 66666
rect 35354 66614 35356 66666
rect 35300 66612 35356 66614
rect 35404 66666 35460 66668
rect 35404 66614 35406 66666
rect 35406 66614 35458 66666
rect 35458 66614 35460 66666
rect 35404 66612 35460 66614
rect 65916 66666 65972 66668
rect 65916 66614 65918 66666
rect 65918 66614 65970 66666
rect 65970 66614 65972 66666
rect 65916 66612 65972 66614
rect 66020 66666 66076 66668
rect 66020 66614 66022 66666
rect 66022 66614 66074 66666
rect 66074 66614 66076 66666
rect 66020 66612 66076 66614
rect 66124 66666 66180 66668
rect 66124 66614 66126 66666
rect 66126 66614 66178 66666
rect 66178 66614 66180 66666
rect 66124 66612 66180 66614
rect 19836 65882 19892 65884
rect 19836 65830 19838 65882
rect 19838 65830 19890 65882
rect 19890 65830 19892 65882
rect 19836 65828 19892 65830
rect 19940 65882 19996 65884
rect 19940 65830 19942 65882
rect 19942 65830 19994 65882
rect 19994 65830 19996 65882
rect 19940 65828 19996 65830
rect 20044 65882 20100 65884
rect 20044 65830 20046 65882
rect 20046 65830 20098 65882
rect 20098 65830 20100 65882
rect 20044 65828 20100 65830
rect 50556 65882 50612 65884
rect 50556 65830 50558 65882
rect 50558 65830 50610 65882
rect 50610 65830 50612 65882
rect 50556 65828 50612 65830
rect 50660 65882 50716 65884
rect 50660 65830 50662 65882
rect 50662 65830 50714 65882
rect 50714 65830 50716 65882
rect 50660 65828 50716 65830
rect 50764 65882 50820 65884
rect 50764 65830 50766 65882
rect 50766 65830 50818 65882
rect 50818 65830 50820 65882
rect 50764 65828 50820 65830
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 35196 65098 35252 65100
rect 35196 65046 35198 65098
rect 35198 65046 35250 65098
rect 35250 65046 35252 65098
rect 35196 65044 35252 65046
rect 35300 65098 35356 65100
rect 35300 65046 35302 65098
rect 35302 65046 35354 65098
rect 35354 65046 35356 65098
rect 35300 65044 35356 65046
rect 35404 65098 35460 65100
rect 35404 65046 35406 65098
rect 35406 65046 35458 65098
rect 35458 65046 35460 65098
rect 35404 65044 35460 65046
rect 65916 65098 65972 65100
rect 65916 65046 65918 65098
rect 65918 65046 65970 65098
rect 65970 65046 65972 65098
rect 65916 65044 65972 65046
rect 66020 65098 66076 65100
rect 66020 65046 66022 65098
rect 66022 65046 66074 65098
rect 66074 65046 66076 65098
rect 66020 65044 66076 65046
rect 66124 65098 66180 65100
rect 66124 65046 66126 65098
rect 66126 65046 66178 65098
rect 66178 65046 66180 65098
rect 66124 65044 66180 65046
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 50556 64314 50612 64316
rect 50556 64262 50558 64314
rect 50558 64262 50610 64314
rect 50610 64262 50612 64314
rect 50556 64260 50612 64262
rect 50660 64314 50716 64316
rect 50660 64262 50662 64314
rect 50662 64262 50714 64314
rect 50714 64262 50716 64314
rect 50660 64260 50716 64262
rect 50764 64314 50820 64316
rect 50764 64262 50766 64314
rect 50766 64262 50818 64314
rect 50818 64262 50820 64314
rect 50764 64260 50820 64262
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 35404 63476 35460 63478
rect 65916 63530 65972 63532
rect 65916 63478 65918 63530
rect 65918 63478 65970 63530
rect 65970 63478 65972 63530
rect 65916 63476 65972 63478
rect 66020 63530 66076 63532
rect 66020 63478 66022 63530
rect 66022 63478 66074 63530
rect 66074 63478 66076 63530
rect 66020 63476 66076 63478
rect 66124 63530 66180 63532
rect 66124 63478 66126 63530
rect 66126 63478 66178 63530
rect 66178 63478 66180 63530
rect 66124 63476 66180 63478
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 50556 62746 50612 62748
rect 50556 62694 50558 62746
rect 50558 62694 50610 62746
rect 50610 62694 50612 62746
rect 50556 62692 50612 62694
rect 50660 62746 50716 62748
rect 50660 62694 50662 62746
rect 50662 62694 50714 62746
rect 50714 62694 50716 62746
rect 50660 62692 50716 62694
rect 50764 62746 50820 62748
rect 50764 62694 50766 62746
rect 50766 62694 50818 62746
rect 50818 62694 50820 62746
rect 50764 62692 50820 62694
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 65916 61962 65972 61964
rect 65916 61910 65918 61962
rect 65918 61910 65970 61962
rect 65970 61910 65972 61962
rect 65916 61908 65972 61910
rect 66020 61962 66076 61964
rect 66020 61910 66022 61962
rect 66022 61910 66074 61962
rect 66074 61910 66076 61962
rect 66020 61908 66076 61910
rect 66124 61962 66180 61964
rect 66124 61910 66126 61962
rect 66126 61910 66178 61962
rect 66178 61910 66180 61962
rect 66124 61908 66180 61910
rect 19836 61178 19892 61180
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 50556 61178 50612 61180
rect 50556 61126 50558 61178
rect 50558 61126 50610 61178
rect 50610 61126 50612 61178
rect 50556 61124 50612 61126
rect 50660 61178 50716 61180
rect 50660 61126 50662 61178
rect 50662 61126 50714 61178
rect 50714 61126 50716 61178
rect 50660 61124 50716 61126
rect 50764 61178 50820 61180
rect 50764 61126 50766 61178
rect 50766 61126 50818 61178
rect 50818 61126 50820 61178
rect 50764 61124 50820 61126
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 65916 60394 65972 60396
rect 65916 60342 65918 60394
rect 65918 60342 65970 60394
rect 65970 60342 65972 60394
rect 65916 60340 65972 60342
rect 66020 60394 66076 60396
rect 66020 60342 66022 60394
rect 66022 60342 66074 60394
rect 66074 60342 66076 60394
rect 66020 60340 66076 60342
rect 66124 60394 66180 60396
rect 66124 60342 66126 60394
rect 66126 60342 66178 60394
rect 66178 60342 66180 60394
rect 66124 60340 66180 60342
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 50556 59610 50612 59612
rect 50556 59558 50558 59610
rect 50558 59558 50610 59610
rect 50610 59558 50612 59610
rect 50556 59556 50612 59558
rect 50660 59610 50716 59612
rect 50660 59558 50662 59610
rect 50662 59558 50714 59610
rect 50714 59558 50716 59610
rect 50660 59556 50716 59558
rect 50764 59610 50820 59612
rect 50764 59558 50766 59610
rect 50766 59558 50818 59610
rect 50818 59558 50820 59610
rect 50764 59556 50820 59558
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 65916 58826 65972 58828
rect 65916 58774 65918 58826
rect 65918 58774 65970 58826
rect 65970 58774 65972 58826
rect 65916 58772 65972 58774
rect 66020 58826 66076 58828
rect 66020 58774 66022 58826
rect 66022 58774 66074 58826
rect 66074 58774 66076 58826
rect 66020 58772 66076 58774
rect 66124 58826 66180 58828
rect 66124 58774 66126 58826
rect 66126 58774 66178 58826
rect 66178 58774 66180 58826
rect 66124 58772 66180 58774
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 50556 58042 50612 58044
rect 50556 57990 50558 58042
rect 50558 57990 50610 58042
rect 50610 57990 50612 58042
rect 50556 57988 50612 57990
rect 50660 58042 50716 58044
rect 50660 57990 50662 58042
rect 50662 57990 50714 58042
rect 50714 57990 50716 58042
rect 50660 57988 50716 57990
rect 50764 58042 50820 58044
rect 50764 57990 50766 58042
rect 50766 57990 50818 58042
rect 50818 57990 50820 58042
rect 50764 57988 50820 57990
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 65916 57258 65972 57260
rect 65916 57206 65918 57258
rect 65918 57206 65970 57258
rect 65970 57206 65972 57258
rect 65916 57204 65972 57206
rect 66020 57258 66076 57260
rect 66020 57206 66022 57258
rect 66022 57206 66074 57258
rect 66074 57206 66076 57258
rect 66020 57204 66076 57206
rect 66124 57258 66180 57260
rect 66124 57206 66126 57258
rect 66126 57206 66178 57258
rect 66178 57206 66180 57258
rect 66124 57204 66180 57206
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 65916 55690 65972 55692
rect 65916 55638 65918 55690
rect 65918 55638 65970 55690
rect 65970 55638 65972 55690
rect 65916 55636 65972 55638
rect 66020 55690 66076 55692
rect 66020 55638 66022 55690
rect 66022 55638 66074 55690
rect 66074 55638 66076 55690
rect 66020 55636 66076 55638
rect 66124 55690 66180 55692
rect 66124 55638 66126 55690
rect 66126 55638 66178 55690
rect 66178 55638 66180 55690
rect 66124 55636 66180 55638
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 65916 54122 65972 54124
rect 65916 54070 65918 54122
rect 65918 54070 65970 54122
rect 65970 54070 65972 54122
rect 65916 54068 65972 54070
rect 66020 54122 66076 54124
rect 66020 54070 66022 54122
rect 66022 54070 66074 54122
rect 66074 54070 66076 54122
rect 66020 54068 66076 54070
rect 66124 54122 66180 54124
rect 66124 54070 66126 54122
rect 66126 54070 66178 54122
rect 66178 54070 66180 54122
rect 66124 54068 66180 54070
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 65916 52554 65972 52556
rect 65916 52502 65918 52554
rect 65918 52502 65970 52554
rect 65970 52502 65972 52554
rect 65916 52500 65972 52502
rect 66020 52554 66076 52556
rect 66020 52502 66022 52554
rect 66022 52502 66074 52554
rect 66074 52502 66076 52554
rect 66020 52500 66076 52502
rect 66124 52554 66180 52556
rect 66124 52502 66126 52554
rect 66126 52502 66178 52554
rect 66178 52502 66180 52554
rect 66124 52500 66180 52502
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 65916 50986 65972 50988
rect 65916 50934 65918 50986
rect 65918 50934 65970 50986
rect 65970 50934 65972 50986
rect 65916 50932 65972 50934
rect 66020 50986 66076 50988
rect 66020 50934 66022 50986
rect 66022 50934 66074 50986
rect 66074 50934 66076 50986
rect 66020 50932 66076 50934
rect 66124 50986 66180 50988
rect 66124 50934 66126 50986
rect 66126 50934 66178 50986
rect 66178 50934 66180 50986
rect 66124 50932 66180 50934
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 65916 49418 65972 49420
rect 65916 49366 65918 49418
rect 65918 49366 65970 49418
rect 65970 49366 65972 49418
rect 65916 49364 65972 49366
rect 66020 49418 66076 49420
rect 66020 49366 66022 49418
rect 66022 49366 66074 49418
rect 66074 49366 66076 49418
rect 66020 49364 66076 49366
rect 66124 49418 66180 49420
rect 66124 49366 66126 49418
rect 66126 49366 66178 49418
rect 66178 49366 66180 49418
rect 66124 49364 66180 49366
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 65916 47850 65972 47852
rect 65916 47798 65918 47850
rect 65918 47798 65970 47850
rect 65970 47798 65972 47850
rect 65916 47796 65972 47798
rect 66020 47850 66076 47852
rect 66020 47798 66022 47850
rect 66022 47798 66074 47850
rect 66074 47798 66076 47850
rect 66020 47796 66076 47798
rect 66124 47850 66180 47852
rect 66124 47798 66126 47850
rect 66126 47798 66178 47850
rect 66178 47798 66180 47850
rect 66124 47796 66180 47798
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 65916 46282 65972 46284
rect 65916 46230 65918 46282
rect 65918 46230 65970 46282
rect 65970 46230 65972 46282
rect 65916 46228 65972 46230
rect 66020 46282 66076 46284
rect 66020 46230 66022 46282
rect 66022 46230 66074 46282
rect 66074 46230 66076 46282
rect 66020 46228 66076 46230
rect 66124 46282 66180 46284
rect 66124 46230 66126 46282
rect 66126 46230 66178 46282
rect 66178 46230 66180 46282
rect 66124 46228 66180 46230
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 65916 44714 65972 44716
rect 65916 44662 65918 44714
rect 65918 44662 65970 44714
rect 65970 44662 65972 44714
rect 65916 44660 65972 44662
rect 66020 44714 66076 44716
rect 66020 44662 66022 44714
rect 66022 44662 66074 44714
rect 66074 44662 66076 44714
rect 66020 44660 66076 44662
rect 66124 44714 66180 44716
rect 66124 44662 66126 44714
rect 66126 44662 66178 44714
rect 66178 44662 66180 44714
rect 66124 44660 66180 44662
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 65916 43146 65972 43148
rect 65916 43094 65918 43146
rect 65918 43094 65970 43146
rect 65970 43094 65972 43146
rect 65916 43092 65972 43094
rect 66020 43146 66076 43148
rect 66020 43094 66022 43146
rect 66022 43094 66074 43146
rect 66074 43094 66076 43146
rect 66020 43092 66076 43094
rect 66124 43146 66180 43148
rect 66124 43094 66126 43146
rect 66126 43094 66178 43146
rect 66178 43094 66180 43146
rect 66124 43092 66180 43094
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 65916 41578 65972 41580
rect 65916 41526 65918 41578
rect 65918 41526 65970 41578
rect 65970 41526 65972 41578
rect 65916 41524 65972 41526
rect 66020 41578 66076 41580
rect 66020 41526 66022 41578
rect 66022 41526 66074 41578
rect 66074 41526 66076 41578
rect 66020 41524 66076 41526
rect 66124 41578 66180 41580
rect 66124 41526 66126 41578
rect 66126 41526 66178 41578
rect 66178 41526 66180 41578
rect 66124 41524 66180 41526
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 65916 40010 65972 40012
rect 65916 39958 65918 40010
rect 65918 39958 65970 40010
rect 65970 39958 65972 40010
rect 65916 39956 65972 39958
rect 66020 40010 66076 40012
rect 66020 39958 66022 40010
rect 66022 39958 66074 40010
rect 66074 39958 66076 40010
rect 66020 39956 66076 39958
rect 66124 40010 66180 40012
rect 66124 39958 66126 40010
rect 66126 39958 66178 40010
rect 66178 39958 66180 40010
rect 66124 39956 66180 39958
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 65916 38442 65972 38444
rect 65916 38390 65918 38442
rect 65918 38390 65970 38442
rect 65970 38390 65972 38442
rect 65916 38388 65972 38390
rect 66020 38442 66076 38444
rect 66020 38390 66022 38442
rect 66022 38390 66074 38442
rect 66074 38390 66076 38442
rect 66020 38388 66076 38390
rect 66124 38442 66180 38444
rect 66124 38390 66126 38442
rect 66126 38390 66178 38442
rect 66178 38390 66180 38442
rect 66124 38388 66180 38390
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 65916 36874 65972 36876
rect 65916 36822 65918 36874
rect 65918 36822 65970 36874
rect 65970 36822 65972 36874
rect 65916 36820 65972 36822
rect 66020 36874 66076 36876
rect 66020 36822 66022 36874
rect 66022 36822 66074 36874
rect 66074 36822 66076 36874
rect 66020 36820 66076 36822
rect 66124 36874 66180 36876
rect 66124 36822 66126 36874
rect 66126 36822 66178 36874
rect 66178 36822 66180 36874
rect 66124 36820 66180 36822
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 65916 35306 65972 35308
rect 65916 35254 65918 35306
rect 65918 35254 65970 35306
rect 65970 35254 65972 35306
rect 65916 35252 65972 35254
rect 66020 35306 66076 35308
rect 66020 35254 66022 35306
rect 66022 35254 66074 35306
rect 66074 35254 66076 35306
rect 66020 35252 66076 35254
rect 66124 35306 66180 35308
rect 66124 35254 66126 35306
rect 66126 35254 66178 35306
rect 66178 35254 66180 35306
rect 66124 35252 66180 35254
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 65916 33738 65972 33740
rect 65916 33686 65918 33738
rect 65918 33686 65970 33738
rect 65970 33686 65972 33738
rect 65916 33684 65972 33686
rect 66020 33738 66076 33740
rect 66020 33686 66022 33738
rect 66022 33686 66074 33738
rect 66074 33686 66076 33738
rect 66020 33684 66076 33686
rect 66124 33738 66180 33740
rect 66124 33686 66126 33738
rect 66126 33686 66178 33738
rect 66178 33686 66180 33738
rect 66124 33684 66180 33686
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 65916 32170 65972 32172
rect 65916 32118 65918 32170
rect 65918 32118 65970 32170
rect 65970 32118 65972 32170
rect 65916 32116 65972 32118
rect 66020 32170 66076 32172
rect 66020 32118 66022 32170
rect 66022 32118 66074 32170
rect 66074 32118 66076 32170
rect 66020 32116 66076 32118
rect 66124 32170 66180 32172
rect 66124 32118 66126 32170
rect 66126 32118 66178 32170
rect 66178 32118 66180 32170
rect 66124 32116 66180 32118
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 65916 30602 65972 30604
rect 65916 30550 65918 30602
rect 65918 30550 65970 30602
rect 65970 30550 65972 30602
rect 65916 30548 65972 30550
rect 66020 30602 66076 30604
rect 66020 30550 66022 30602
rect 66022 30550 66074 30602
rect 66074 30550 66076 30602
rect 66020 30548 66076 30550
rect 66124 30602 66180 30604
rect 66124 30550 66126 30602
rect 66126 30550 66178 30602
rect 66178 30550 66180 30602
rect 66124 30548 66180 30550
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 65916 29034 65972 29036
rect 65916 28982 65918 29034
rect 65918 28982 65970 29034
rect 65970 28982 65972 29034
rect 65916 28980 65972 28982
rect 66020 29034 66076 29036
rect 66020 28982 66022 29034
rect 66022 28982 66074 29034
rect 66074 28982 66076 29034
rect 66020 28980 66076 28982
rect 66124 29034 66180 29036
rect 66124 28982 66126 29034
rect 66126 28982 66178 29034
rect 66178 28982 66180 29034
rect 66124 28980 66180 28982
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 65916 27466 65972 27468
rect 65916 27414 65918 27466
rect 65918 27414 65970 27466
rect 65970 27414 65972 27466
rect 65916 27412 65972 27414
rect 66020 27466 66076 27468
rect 66020 27414 66022 27466
rect 66022 27414 66074 27466
rect 66074 27414 66076 27466
rect 66020 27412 66076 27414
rect 66124 27466 66180 27468
rect 66124 27414 66126 27466
rect 66126 27414 66178 27466
rect 66178 27414 66180 27466
rect 66124 27412 66180 27414
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 65916 25898 65972 25900
rect 65916 25846 65918 25898
rect 65918 25846 65970 25898
rect 65970 25846 65972 25898
rect 65916 25844 65972 25846
rect 66020 25898 66076 25900
rect 66020 25846 66022 25898
rect 66022 25846 66074 25898
rect 66074 25846 66076 25898
rect 66020 25844 66076 25846
rect 66124 25898 66180 25900
rect 66124 25846 66126 25898
rect 66126 25846 66178 25898
rect 66178 25846 66180 25898
rect 66124 25844 66180 25846
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 65916 24330 65972 24332
rect 65916 24278 65918 24330
rect 65918 24278 65970 24330
rect 65970 24278 65972 24330
rect 65916 24276 65972 24278
rect 66020 24330 66076 24332
rect 66020 24278 66022 24330
rect 66022 24278 66074 24330
rect 66074 24278 66076 24330
rect 66020 24276 66076 24278
rect 66124 24330 66180 24332
rect 66124 24278 66126 24330
rect 66126 24278 66178 24330
rect 66178 24278 66180 24330
rect 66124 24276 66180 24278
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 65916 22762 65972 22764
rect 65916 22710 65918 22762
rect 65918 22710 65970 22762
rect 65970 22710 65972 22762
rect 65916 22708 65972 22710
rect 66020 22762 66076 22764
rect 66020 22710 66022 22762
rect 66022 22710 66074 22762
rect 66074 22710 66076 22762
rect 66020 22708 66076 22710
rect 66124 22762 66180 22764
rect 66124 22710 66126 22762
rect 66126 22710 66178 22762
rect 66178 22710 66180 22762
rect 66124 22708 66180 22710
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 65916 21194 65972 21196
rect 65916 21142 65918 21194
rect 65918 21142 65970 21194
rect 65970 21142 65972 21194
rect 65916 21140 65972 21142
rect 66020 21194 66076 21196
rect 66020 21142 66022 21194
rect 66022 21142 66074 21194
rect 66074 21142 66076 21194
rect 66020 21140 66076 21142
rect 66124 21194 66180 21196
rect 66124 21142 66126 21194
rect 66126 21142 66178 21194
rect 66178 21142 66180 21194
rect 66124 21140 66180 21142
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 65916 19626 65972 19628
rect 65916 19574 65918 19626
rect 65918 19574 65970 19626
rect 65970 19574 65972 19626
rect 65916 19572 65972 19574
rect 66020 19626 66076 19628
rect 66020 19574 66022 19626
rect 66022 19574 66074 19626
rect 66074 19574 66076 19626
rect 66020 19572 66076 19574
rect 66124 19626 66180 19628
rect 66124 19574 66126 19626
rect 66126 19574 66178 19626
rect 66178 19574 66180 19626
rect 66124 19572 66180 19574
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 65916 18058 65972 18060
rect 65916 18006 65918 18058
rect 65918 18006 65970 18058
rect 65970 18006 65972 18058
rect 65916 18004 65972 18006
rect 66020 18058 66076 18060
rect 66020 18006 66022 18058
rect 66022 18006 66074 18058
rect 66074 18006 66076 18058
rect 66020 18004 66076 18006
rect 66124 18058 66180 18060
rect 66124 18006 66126 18058
rect 66126 18006 66178 18058
rect 66178 18006 66180 18058
rect 66124 18004 66180 18006
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 65916 16490 65972 16492
rect 65916 16438 65918 16490
rect 65918 16438 65970 16490
rect 65970 16438 65972 16490
rect 65916 16436 65972 16438
rect 66020 16490 66076 16492
rect 66020 16438 66022 16490
rect 66022 16438 66074 16490
rect 66074 16438 66076 16490
rect 66020 16436 66076 16438
rect 66124 16490 66180 16492
rect 66124 16438 66126 16490
rect 66126 16438 66178 16490
rect 66178 16438 66180 16490
rect 66124 16436 66180 16438
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 65916 14922 65972 14924
rect 65916 14870 65918 14922
rect 65918 14870 65970 14922
rect 65970 14870 65972 14922
rect 65916 14868 65972 14870
rect 66020 14922 66076 14924
rect 66020 14870 66022 14922
rect 66022 14870 66074 14922
rect 66074 14870 66076 14922
rect 66020 14868 66076 14870
rect 66124 14922 66180 14924
rect 66124 14870 66126 14922
rect 66126 14870 66178 14922
rect 66178 14870 66180 14922
rect 66124 14868 66180 14870
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 65916 13354 65972 13356
rect 65916 13302 65918 13354
rect 65918 13302 65970 13354
rect 65970 13302 65972 13354
rect 65916 13300 65972 13302
rect 66020 13354 66076 13356
rect 66020 13302 66022 13354
rect 66022 13302 66074 13354
rect 66074 13302 66076 13354
rect 66020 13300 66076 13302
rect 66124 13354 66180 13356
rect 66124 13302 66126 13354
rect 66126 13302 66178 13354
rect 66178 13302 66180 13354
rect 66124 13300 66180 13302
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 65916 11786 65972 11788
rect 65916 11734 65918 11786
rect 65918 11734 65970 11786
rect 65970 11734 65972 11786
rect 65916 11732 65972 11734
rect 66020 11786 66076 11788
rect 66020 11734 66022 11786
rect 66022 11734 66074 11786
rect 66074 11734 66076 11786
rect 66020 11732 66076 11734
rect 66124 11786 66180 11788
rect 66124 11734 66126 11786
rect 66126 11734 66178 11786
rect 66178 11734 66180 11786
rect 66124 11732 66180 11734
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 65916 10218 65972 10220
rect 65916 10166 65918 10218
rect 65918 10166 65970 10218
rect 65970 10166 65972 10218
rect 65916 10164 65972 10166
rect 66020 10218 66076 10220
rect 66020 10166 66022 10218
rect 66022 10166 66074 10218
rect 66074 10166 66076 10218
rect 66020 10164 66076 10166
rect 66124 10218 66180 10220
rect 66124 10166 66126 10218
rect 66126 10166 66178 10218
rect 66178 10166 66180 10218
rect 66124 10164 66180 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 65916 8650 65972 8652
rect 65916 8598 65918 8650
rect 65918 8598 65970 8650
rect 65970 8598 65972 8650
rect 65916 8596 65972 8598
rect 66020 8650 66076 8652
rect 66020 8598 66022 8650
rect 66022 8598 66074 8650
rect 66074 8598 66076 8650
rect 66020 8596 66076 8598
rect 66124 8650 66180 8652
rect 66124 8598 66126 8650
rect 66126 8598 66178 8650
rect 66178 8598 66180 8650
rect 66124 8596 66180 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 65916 7082 65972 7084
rect 65916 7030 65918 7082
rect 65918 7030 65970 7082
rect 65970 7030 65972 7082
rect 65916 7028 65972 7030
rect 66020 7082 66076 7084
rect 66020 7030 66022 7082
rect 66022 7030 66074 7082
rect 66074 7030 66076 7082
rect 66020 7028 66076 7030
rect 66124 7082 66180 7084
rect 66124 7030 66126 7082
rect 66126 7030 66178 7082
rect 66178 7030 66180 7082
rect 66124 7028 66180 7030
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 65916 5514 65972 5516
rect 65916 5462 65918 5514
rect 65918 5462 65970 5514
rect 65970 5462 65972 5514
rect 65916 5460 65972 5462
rect 66020 5514 66076 5516
rect 66020 5462 66022 5514
rect 66022 5462 66074 5514
rect 66074 5462 66076 5514
rect 66020 5460 66076 5462
rect 66124 5514 66180 5516
rect 66124 5462 66126 5514
rect 66126 5462 66178 5514
rect 66178 5462 66180 5514
rect 66124 5460 66180 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 65916 3946 65972 3948
rect 65916 3894 65918 3946
rect 65918 3894 65970 3946
rect 65970 3894 65972 3946
rect 65916 3892 65972 3894
rect 66020 3946 66076 3948
rect 66020 3894 66022 3946
rect 66022 3894 66074 3946
rect 66074 3894 66076 3946
rect 66020 3892 66076 3894
rect 66124 3946 66180 3948
rect 66124 3894 66126 3946
rect 66126 3894 66178 3946
rect 66178 3894 66180 3946
rect 66124 3892 66180 3894
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 41804 3276 41860 3332
rect 42364 3330 42420 3332
rect 42364 3278 42366 3330
rect 42366 3278 42418 3330
rect 42418 3278 42420 3330
rect 42364 3276 42420 3278
rect 43148 3276 43204 3332
rect 43708 3330 43764 3332
rect 43708 3278 43710 3330
rect 43710 3278 43762 3330
rect 43762 3278 43764 3330
rect 43708 3276 43764 3278
rect 45164 3276 45220 3332
rect 45724 3330 45780 3332
rect 45724 3278 45726 3330
rect 45726 3278 45778 3330
rect 45778 3278 45780 3330
rect 45724 3276 45780 3278
rect 46508 3276 46564 3332
rect 47068 3330 47124 3332
rect 47068 3278 47070 3330
rect 47070 3278 47122 3330
rect 47122 3278 47124 3330
rect 47068 3276 47124 3278
rect 48524 3276 48580 3332
rect 49084 3330 49140 3332
rect 49084 3278 49086 3330
rect 49086 3278 49138 3330
rect 49138 3278 49140 3330
rect 49084 3276 49140 3278
rect 49868 3276 49924 3332
rect 50428 3330 50484 3332
rect 50428 3278 50430 3330
rect 50430 3278 50482 3330
rect 50482 3278 50484 3330
rect 50428 3276 50484 3278
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 51884 3276 51940 3332
rect 52444 3330 52500 3332
rect 52444 3278 52446 3330
rect 52446 3278 52498 3330
rect 52498 3278 52500 3330
rect 52444 3276 52500 3278
rect 53228 3276 53284 3332
rect 53788 3330 53844 3332
rect 53788 3278 53790 3330
rect 53790 3278 53842 3330
rect 53842 3278 53844 3330
rect 53788 3276 53844 3278
rect 55132 1708 55188 1764
rect 55804 1708 55860 1764
rect 56588 3276 56644 3332
rect 57148 3330 57204 3332
rect 57148 3278 57150 3330
rect 57150 3278 57202 3330
rect 57202 3278 57204 3330
rect 57148 3276 57204 3278
rect 58604 3276 58660 3332
rect 59164 3330 59220 3332
rect 59164 3278 59166 3330
rect 59166 3278 59218 3330
rect 59218 3278 59220 3330
rect 59164 3276 59220 3278
rect 59948 3276 60004 3332
rect 60508 3330 60564 3332
rect 60508 3278 60510 3330
rect 60510 3278 60562 3330
rect 60562 3278 60564 3330
rect 60508 3276 60564 3278
rect 61180 3276 61236 3332
rect 62300 3330 62356 3332
rect 62300 3278 62302 3330
rect 62302 3278 62354 3330
rect 62354 3278 62356 3330
rect 62300 3276 62356 3278
rect 61852 1708 61908 1764
rect 62972 1708 63028 1764
rect 63196 3276 63252 3332
rect 64316 3330 64372 3332
rect 64316 3278 64318 3330
rect 64318 3278 64370 3330
rect 64370 3278 64372 3330
rect 64316 3276 64372 3278
rect 64540 3276 64596 3332
rect 65660 3330 65716 3332
rect 65660 3278 65662 3330
rect 65662 3278 65714 3330
rect 65714 3278 65716 3330
rect 65660 3276 65716 3278
rect 65212 1708 65268 1764
rect 66332 1708 66388 1764
rect 66556 3276 66612 3332
rect 67676 3330 67732 3332
rect 67676 3278 67678 3330
rect 67678 3278 67730 3330
rect 67730 3278 67732 3330
rect 67676 3276 67732 3278
rect 67900 3276 67956 3332
rect 69020 3330 69076 3332
rect 69020 3278 69022 3330
rect 69022 3278 69074 3330
rect 69074 3278 69076 3330
rect 69020 3276 69076 3278
rect 68572 1708 68628 1764
rect 69692 1708 69748 1764
rect 69916 3276 69972 3332
rect 71036 3330 71092 3332
rect 71036 3278 71038 3330
rect 71038 3278 71090 3330
rect 71090 3278 71092 3330
rect 71036 3276 71092 3278
rect 71260 3276 71316 3332
rect 72380 3330 72436 3332
rect 72380 3278 72382 3330
rect 72382 3278 72434 3330
rect 72434 3278 72436 3330
rect 72380 3276 72436 3278
rect 71932 1708 71988 1764
rect 73052 1708 73108 1764
rect 73388 3276 73444 3332
rect 74396 3330 74452 3332
rect 74396 3278 74398 3330
rect 74398 3278 74450 3330
rect 74450 3278 74452 3330
rect 74396 3276 74452 3278
<< metal3 >>
rect 33170 77532 33180 77588
rect 33236 77532 56588 77588
rect 56644 77532 56654 77588
rect 45826 77420 45836 77476
rect 45892 77420 46956 77476
rect 47012 77420 70924 77476
rect 70980 77420 70990 77476
rect 6514 77308 6524 77364
rect 6580 77308 43708 77364
rect 43764 77308 43774 77364
rect 54002 77308 54012 77364
rect 54068 77308 60620 77364
rect 60676 77308 60686 77364
rect 35746 77196 35756 77252
rect 35812 77196 53228 77252
rect 53284 77196 53294 77252
rect 50642 76972 50652 77028
rect 50708 76972 51548 77028
rect 51604 76972 52892 77028
rect 52948 76972 52958 77028
rect 19826 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20110 76860
rect 50546 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50830 76860
rect 37874 76748 37884 76804
rect 37940 76748 38780 76804
rect 38836 76748 38846 76804
rect 68786 76748 68796 76804
rect 68852 76748 69356 76804
rect 69412 76748 70476 76804
rect 70532 76748 70542 76804
rect 38322 76636 38332 76692
rect 38388 76636 43820 76692
rect 43876 76636 43886 76692
rect 53330 76636 53340 76692
rect 53396 76636 60508 76692
rect 60564 76636 60574 76692
rect 68114 76636 68124 76692
rect 68180 76636 69916 76692
rect 69972 76636 69982 76692
rect 26786 76524 26796 76580
rect 26852 76524 27244 76580
rect 27300 76524 33068 76580
rect 33124 76524 33134 76580
rect 38546 76524 38556 76580
rect 38612 76524 39116 76580
rect 39172 76524 39182 76580
rect 45042 76524 45052 76580
rect 45108 76524 45500 76580
rect 45556 76524 45566 76580
rect 48514 76524 48524 76580
rect 48580 76524 53900 76580
rect 53956 76524 53966 76580
rect 56690 76524 56700 76580
rect 56756 76524 57932 76580
rect 57988 76524 58604 76580
rect 58660 76524 58670 76580
rect 62738 76524 62748 76580
rect 62804 76524 63532 76580
rect 63588 76524 64988 76580
rect 65044 76524 65054 76580
rect 65202 76524 65212 76580
rect 65268 76524 68012 76580
rect 68068 76524 68078 76580
rect 70802 76524 70812 76580
rect 70868 76524 73052 76580
rect 73108 76524 73118 76580
rect 5058 76412 5068 76468
rect 5124 76412 6524 76468
rect 6580 76412 6590 76468
rect 13122 76412 13132 76468
rect 13188 76412 13804 76468
rect 13860 76412 13870 76468
rect 15138 76412 15148 76468
rect 15204 76412 15820 76468
rect 15876 76412 15886 76468
rect 24994 76412 25004 76468
rect 25060 76412 29260 76468
rect 29316 76412 29326 76468
rect 34626 76412 34636 76468
rect 34692 76412 36092 76468
rect 36148 76412 36158 76468
rect 45938 76412 45948 76468
rect 46004 76412 46956 76468
rect 47012 76412 47022 76468
rect 51986 76412 51996 76468
rect 52052 76412 59836 76468
rect 59892 76412 59902 76468
rect 60060 76412 62412 76468
rect 62468 76412 62478 76468
rect 60060 76356 60116 76412
rect 27794 76300 27804 76356
rect 27860 76300 28812 76356
rect 28868 76300 28878 76356
rect 29810 76300 29820 76356
rect 29876 76300 30716 76356
rect 30772 76300 30782 76356
rect 31826 76300 31836 76356
rect 31892 76300 32732 76356
rect 32788 76300 32798 76356
rect 39330 76300 39340 76356
rect 39396 76300 41692 76356
rect 41748 76300 41758 76356
rect 42802 76300 42812 76356
rect 42868 76300 46396 76356
rect 46452 76300 49084 76356
rect 49140 76300 49150 76356
rect 52658 76300 52668 76356
rect 52724 76300 54236 76356
rect 54292 76300 60116 76356
rect 60274 76300 60284 76356
rect 60340 76300 69020 76356
rect 69076 76300 69086 76356
rect 20962 76188 20972 76244
rect 21028 76188 35084 76244
rect 35140 76188 35150 76244
rect 35970 76188 35980 76244
rect 36036 76188 40012 76244
rect 40068 76188 44044 76244
rect 44100 76188 44716 76244
rect 44772 76188 44782 76244
rect 60396 76188 62860 76244
rect 62916 76188 62926 76244
rect 63084 76188 74508 76244
rect 74564 76188 74574 76244
rect 23202 76076 23212 76132
rect 23268 76076 23996 76132
rect 24052 76076 34356 76132
rect 36642 76076 36652 76132
rect 36708 76076 48972 76132
rect 49028 76076 49038 76132
rect 58370 76076 58380 76132
rect 58436 76076 60172 76132
rect 60228 76076 60238 76132
rect 4466 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4750 76076
rect 29474 75964 29484 76020
rect 29540 75964 32172 76020
rect 32228 75964 32238 76020
rect 34300 75908 34356 76076
rect 35186 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35470 76076
rect 37986 75964 37996 76020
rect 38052 75964 45500 76020
rect 45556 75964 48412 76020
rect 48468 75964 48478 76020
rect 52322 75964 52332 76020
rect 52388 75964 54348 76020
rect 54404 75964 59612 76020
rect 59668 75964 59678 76020
rect 60396 75908 60452 76188
rect 63084 76132 63140 76188
rect 62514 76076 62524 76132
rect 62580 76076 63140 76132
rect 65906 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66190 76076
rect 3378 75852 3388 75908
rect 3444 75852 21644 75908
rect 21700 75852 21710 75908
rect 34300 75852 36316 75908
rect 36372 75852 36382 75908
rect 38882 75852 38892 75908
rect 38948 75852 40236 75908
rect 40292 75852 45052 75908
rect 45108 75852 45118 75908
rect 53106 75852 53116 75908
rect 53172 75852 56140 75908
rect 56196 75852 56206 75908
rect 56354 75852 56364 75908
rect 56420 75852 56924 75908
rect 56980 75852 56990 75908
rect 59154 75852 59164 75908
rect 59220 75852 60452 75908
rect 19170 75740 19180 75796
rect 19236 75740 19852 75796
rect 19908 75740 19918 75796
rect 29362 75740 29372 75796
rect 29428 75740 30828 75796
rect 30884 75740 30894 75796
rect 39862 75740 39900 75796
rect 39956 75740 39966 75796
rect 40450 75740 40460 75796
rect 40516 75740 44828 75796
rect 44884 75740 44894 75796
rect 49074 75740 49084 75796
rect 49140 75740 51100 75796
rect 51156 75740 51166 75796
rect 53554 75740 53564 75796
rect 53620 75740 58940 75796
rect 58996 75740 59006 75796
rect 16930 75628 16940 75684
rect 16996 75628 17836 75684
rect 17892 75628 23492 75684
rect 30034 75628 30044 75684
rect 30100 75628 30492 75684
rect 30548 75628 30558 75684
rect 38658 75628 38668 75684
rect 38724 75628 41132 75684
rect 41188 75628 41198 75684
rect 43922 75628 43932 75684
rect 43988 75628 43998 75684
rect 52994 75628 53004 75684
rect 53060 75628 54124 75684
rect 54180 75628 54190 75684
rect 54450 75628 54460 75684
rect 54516 75628 55132 75684
rect 55188 75628 55198 75684
rect 55346 75628 55356 75684
rect 55412 75628 61628 75684
rect 61684 75628 61694 75684
rect 66556 75628 75068 75684
rect 75124 75628 75134 75684
rect 21074 75516 21084 75572
rect 21140 75516 21756 75572
rect 21812 75516 21822 75572
rect 23436 75460 23492 75628
rect 30258 75516 30268 75572
rect 30324 75516 30604 75572
rect 30660 75516 31164 75572
rect 31220 75516 32060 75572
rect 32116 75516 32126 75572
rect 32610 75516 32620 75572
rect 32676 75516 33852 75572
rect 33908 75516 34076 75572
rect 34132 75516 34142 75572
rect 34402 75516 34412 75572
rect 34468 75516 39900 75572
rect 39956 75516 39966 75572
rect 40450 75516 40460 75572
rect 40516 75516 41692 75572
rect 41748 75516 41758 75572
rect 43026 75516 43036 75572
rect 43092 75516 43260 75572
rect 43316 75516 43484 75572
rect 43540 75516 43550 75572
rect 23436 75404 31276 75460
rect 31332 75404 31342 75460
rect 32274 75404 32284 75460
rect 32340 75404 33180 75460
rect 33236 75404 33246 75460
rect 34290 75404 34300 75460
rect 34356 75404 34972 75460
rect 35028 75404 35756 75460
rect 35812 75404 35822 75460
rect 37538 75404 37548 75460
rect 37604 75404 38612 75460
rect 38668 75404 38678 75460
rect 38770 75404 38780 75460
rect 38836 75404 41244 75460
rect 41300 75404 41310 75460
rect 43670 75404 43708 75460
rect 43764 75404 43774 75460
rect 43932 75348 43988 75628
rect 66556 75572 66612 75628
rect 44482 75516 44492 75572
rect 44548 75516 47404 75572
rect 47460 75516 47470 75572
rect 53778 75516 53788 75572
rect 53844 75516 55580 75572
rect 55636 75516 55646 75572
rect 56466 75516 56476 75572
rect 56532 75516 59948 75572
rect 60004 75516 60014 75572
rect 61394 75516 61404 75572
rect 61460 75516 63084 75572
rect 63140 75516 63150 75572
rect 63858 75516 63868 75572
rect 63924 75516 66612 75572
rect 66770 75516 66780 75572
rect 66836 75516 69020 75572
rect 69076 75516 69086 75572
rect 70130 75516 70140 75572
rect 70196 75516 70700 75572
rect 70756 75516 70766 75572
rect 73490 75516 73500 75572
rect 73556 75516 73948 75572
rect 74004 75516 74014 75572
rect 74946 75516 74956 75572
rect 75012 75516 76972 75572
rect 77028 75516 77420 75572
rect 77476 75516 77486 75572
rect 44146 75404 44156 75460
rect 44212 75404 45612 75460
rect 45668 75404 45678 75460
rect 45938 75404 45948 75460
rect 46004 75404 47180 75460
rect 47236 75404 48300 75460
rect 48356 75404 48366 75460
rect 49074 75404 49084 75460
rect 49140 75404 49756 75460
rect 49812 75404 49822 75460
rect 54002 75404 54012 75460
rect 54068 75404 55020 75460
rect 55076 75404 56140 75460
rect 56196 75404 56206 75460
rect 58034 75404 58044 75460
rect 58100 75404 62412 75460
rect 62468 75404 62478 75460
rect 69458 75404 69468 75460
rect 69524 75404 70028 75460
rect 70084 75404 70094 75460
rect 72818 75404 72828 75460
rect 72884 75404 73388 75460
rect 73444 75404 73454 75460
rect 31892 75292 40124 75348
rect 40180 75292 40190 75348
rect 41122 75292 41132 75348
rect 41188 75292 43596 75348
rect 43652 75292 43662 75348
rect 43932 75292 47404 75348
rect 47460 75292 47470 75348
rect 56018 75292 56028 75348
rect 56084 75292 61740 75348
rect 61796 75292 61806 75348
rect 19826 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20110 75292
rect 31378 75180 31388 75236
rect 31444 75180 31836 75236
rect 31892 75180 31948 75292
rect 50546 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50830 75292
rect 32498 75180 32508 75236
rect 32564 75180 33180 75236
rect 33236 75180 33246 75236
rect 37538 75180 37548 75236
rect 37604 75180 37884 75236
rect 37940 75180 38780 75236
rect 38836 75180 38846 75236
rect 39004 75180 41916 75236
rect 41972 75180 41982 75236
rect 42466 75180 42476 75236
rect 42532 75180 42924 75236
rect 42980 75180 42990 75236
rect 43698 75180 43708 75236
rect 43764 75180 44268 75236
rect 44324 75180 44604 75236
rect 44660 75180 44670 75236
rect 44818 75180 44828 75236
rect 44884 75180 46508 75236
rect 46564 75180 46574 75236
rect 51650 75180 51660 75236
rect 51716 75180 54796 75236
rect 54852 75180 55020 75236
rect 55076 75180 55086 75236
rect 55234 75180 55244 75236
rect 55300 75180 55804 75236
rect 55860 75180 57036 75236
rect 57092 75180 57102 75236
rect 57362 75180 57372 75236
rect 57428 75180 58044 75236
rect 58100 75180 59836 75236
rect 59892 75180 59902 75236
rect 60162 75180 60172 75236
rect 60228 75180 62188 75236
rect 62244 75180 62254 75236
rect 39004 75124 39060 75180
rect 42476 75124 42532 75180
rect 59836 75124 59892 75180
rect 20178 75068 20188 75124
rect 20244 75068 33292 75124
rect 33348 75068 33358 75124
rect 38658 75068 38668 75124
rect 38724 75068 39060 75124
rect 40002 75068 40012 75124
rect 40068 75068 40684 75124
rect 40740 75068 40750 75124
rect 41010 75068 41020 75124
rect 41076 75068 42532 75124
rect 43138 75068 43148 75124
rect 43204 75068 43932 75124
rect 43988 75068 43998 75124
rect 48738 75068 48748 75124
rect 48804 75068 50316 75124
rect 50372 75068 50988 75124
rect 51044 75068 51054 75124
rect 55234 75068 55244 75124
rect 55300 75068 55356 75124
rect 55412 75068 55422 75124
rect 58044 75068 58940 75124
rect 58996 75068 59780 75124
rect 59836 75068 61628 75124
rect 61684 75068 61694 75124
rect 62066 75068 62076 75124
rect 62132 75068 62860 75124
rect 62916 75068 62926 75124
rect 21634 74956 21644 75012
rect 21700 74956 29932 75012
rect 29988 74956 31164 75012
rect 31220 74956 31230 75012
rect 31892 74956 36540 75012
rect 36596 74956 36606 75012
rect 37314 74956 37324 75012
rect 37380 74956 38556 75012
rect 38612 74956 39004 75012
rect 39060 74956 39070 75012
rect 40226 74956 40236 75012
rect 40292 74956 40796 75012
rect 40852 74956 44156 75012
rect 44212 74956 44222 75012
rect 48626 74956 48636 75012
rect 48692 74956 49532 75012
rect 49588 74956 49598 75012
rect 49746 74956 49756 75012
rect 49812 74956 50764 75012
rect 50820 74956 50830 75012
rect 52994 74956 53004 75012
rect 53060 74956 54012 75012
rect 54068 74956 54078 75012
rect 29372 74900 29428 74956
rect 29362 74844 29372 74900
rect 29428 74844 29438 74900
rect 31892 74788 31948 74956
rect 49532 74900 49588 74956
rect 32050 74844 32060 74900
rect 32116 74844 33740 74900
rect 33796 74844 33806 74900
rect 35186 74844 35196 74900
rect 35252 74844 35644 74900
rect 35700 74844 38220 74900
rect 38276 74844 38286 74900
rect 40898 74844 40908 74900
rect 40964 74844 42252 74900
rect 42308 74844 42700 74900
rect 42756 74844 42766 74900
rect 43698 74844 43708 74900
rect 43764 74844 45220 74900
rect 45714 74844 45724 74900
rect 45780 74844 46284 74900
rect 46340 74844 46350 74900
rect 49532 74844 50316 74900
rect 50372 74844 50382 74900
rect 50866 74844 50876 74900
rect 50932 74844 51436 74900
rect 51492 74844 51996 74900
rect 52052 74844 52062 74900
rect 54338 74844 54348 74900
rect 54404 74844 55692 74900
rect 55748 74844 55758 74900
rect 45164 74788 45220 74844
rect 58044 74788 58100 75068
rect 59724 75012 59780 75068
rect 58258 74956 58268 75012
rect 58324 74956 58828 75012
rect 58884 74956 58894 75012
rect 59714 74956 59724 75012
rect 59780 74956 59790 75012
rect 59938 74956 59948 75012
rect 60004 74956 60172 75012
rect 60228 74956 60238 75012
rect 61842 74956 61852 75012
rect 61908 74956 63868 75012
rect 63924 74956 63934 75012
rect 59154 74844 59164 74900
rect 59220 74844 61516 74900
rect 61572 74844 61582 74900
rect 28914 74732 28924 74788
rect 28980 74732 29260 74788
rect 29316 74732 31948 74788
rect 32246 74732 32284 74788
rect 32340 74732 32350 74788
rect 35522 74732 35532 74788
rect 35588 74732 36708 74788
rect 36866 74732 36876 74788
rect 36932 74732 38668 74788
rect 38724 74732 38734 74788
rect 43138 74732 43148 74788
rect 43204 74732 43820 74788
rect 43876 74732 43886 74788
rect 45154 74732 45164 74788
rect 45220 74732 49756 74788
rect 49812 74732 49822 74788
rect 51510 74732 51548 74788
rect 51604 74732 51614 74788
rect 55468 74732 58100 74788
rect 58818 74732 58828 74788
rect 58884 74732 60284 74788
rect 60340 74732 61404 74788
rect 61460 74732 61470 74788
rect 62132 74732 63420 74788
rect 63476 74732 63486 74788
rect 36652 74676 36708 74732
rect 55468 74676 55524 74732
rect 33506 74620 33516 74676
rect 33572 74620 36316 74676
rect 36372 74620 36382 74676
rect 36652 74620 42028 74676
rect 42084 74620 42094 74676
rect 43698 74620 43708 74676
rect 43764 74620 44380 74676
rect 44436 74620 44446 74676
rect 45490 74620 45500 74676
rect 45556 74620 46396 74676
rect 46452 74620 46462 74676
rect 52882 74620 52892 74676
rect 52948 74620 55468 74676
rect 55524 74620 55534 74676
rect 57026 74620 57036 74676
rect 57092 74620 60844 74676
rect 60900 74620 60910 74676
rect 62132 74564 62188 74732
rect 44380 74508 44828 74564
rect 44884 74508 44894 74564
rect 51986 74508 51996 74564
rect 52052 74508 58268 74564
rect 58324 74508 58334 74564
rect 59714 74508 59724 74564
rect 59780 74508 60956 74564
rect 61012 74508 62188 74564
rect 4466 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4750 74508
rect 35186 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35470 74508
rect 44380 74452 44436 74508
rect 65906 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66190 74508
rect 35746 74396 35756 74452
rect 35812 74396 38108 74452
rect 38164 74396 38174 74452
rect 43484 74396 44380 74452
rect 44436 74396 44446 74452
rect 43484 74340 43540 74396
rect 28578 74284 28588 74340
rect 28644 74284 33964 74340
rect 34020 74284 34030 74340
rect 34402 74284 34412 74340
rect 34468 74284 35084 74340
rect 35140 74284 35150 74340
rect 38612 74284 43484 74340
rect 43540 74284 43550 74340
rect 44034 74284 44044 74340
rect 44100 74284 49308 74340
rect 49364 74284 49374 74340
rect 51090 74284 51100 74340
rect 51156 74284 52108 74340
rect 52164 74284 53788 74340
rect 53844 74284 54572 74340
rect 54628 74284 54638 74340
rect 55682 74284 55692 74340
rect 55748 74284 55758 74340
rect 59490 74284 59500 74340
rect 59556 74284 60620 74340
rect 60676 74284 61628 74340
rect 61684 74284 65772 74340
rect 65828 74284 65838 74340
rect 29810 74172 29820 74228
rect 29876 74172 31052 74228
rect 31108 74172 31836 74228
rect 31892 74172 31902 74228
rect 34514 74172 34524 74228
rect 34580 74172 35644 74228
rect 35700 74172 35710 74228
rect 36866 74172 36876 74228
rect 36932 74172 36942 74228
rect 36876 74116 36932 74172
rect 38612 74116 38668 74284
rect 55692 74228 55748 74284
rect 40002 74172 40012 74228
rect 40068 74172 40348 74228
rect 40404 74172 43596 74228
rect 43652 74172 43932 74228
rect 43988 74172 44828 74228
rect 44884 74172 47852 74228
rect 47908 74172 47918 74228
rect 50082 74172 50092 74228
rect 50148 74172 51324 74228
rect 51380 74172 52780 74228
rect 52836 74172 53676 74228
rect 53732 74172 53742 74228
rect 55692 74172 56588 74228
rect 56644 74172 59164 74228
rect 59220 74172 59230 74228
rect 61954 74172 61964 74228
rect 62020 74172 62972 74228
rect 63028 74172 63038 74228
rect 77634 74172 77644 74228
rect 77700 74172 78092 74228
rect 78148 74172 78158 74228
rect 32722 74060 32732 74116
rect 32788 74060 33404 74116
rect 33460 74060 33470 74116
rect 35298 74060 35308 74116
rect 35364 74060 36932 74116
rect 38098 74060 38108 74116
rect 38164 74060 38668 74116
rect 42130 74060 42140 74116
rect 42196 74060 42476 74116
rect 42532 74060 44156 74116
rect 44212 74060 44222 74116
rect 47282 74060 47292 74116
rect 47348 74060 48524 74116
rect 48580 74060 48590 74116
rect 49746 74060 49756 74116
rect 49812 74060 50652 74116
rect 50708 74060 50718 74116
rect 50978 74060 50988 74116
rect 51044 74060 51212 74116
rect 51268 74060 51278 74116
rect 51426 74060 51436 74116
rect 51492 74060 51548 74116
rect 51604 74060 51614 74116
rect 51874 74060 51884 74116
rect 51940 74060 54684 74116
rect 54740 74060 54750 74116
rect 56914 74060 56924 74116
rect 56980 74060 57596 74116
rect 57652 74060 57662 74116
rect 61394 74060 61404 74116
rect 61460 74060 62076 74116
rect 62132 74060 62142 74116
rect 36306 73948 36316 74004
rect 36372 73948 39452 74004
rect 39508 73948 39518 74004
rect 39890 73948 39900 74004
rect 39956 73948 40796 74004
rect 40852 73948 41020 74004
rect 41076 73948 41086 74004
rect 42802 73948 42812 74004
rect 42868 73948 43484 74004
rect 43540 73948 43550 74004
rect 44594 73948 44604 74004
rect 44660 73948 45612 74004
rect 45668 73948 45678 74004
rect 47058 73948 47068 74004
rect 47124 73948 47852 74004
rect 47908 73948 47918 74004
rect 49858 73948 49868 74004
rect 49924 73948 50316 74004
rect 50372 73948 50876 74004
rect 50932 73948 50942 74004
rect 51090 73948 51100 74004
rect 51156 73948 51194 74004
rect 56018 73948 56028 74004
rect 56084 73948 57932 74004
rect 57988 73948 57998 74004
rect 29138 73836 29148 73892
rect 29204 73836 30268 73892
rect 30324 73836 30334 73892
rect 31490 73836 31500 73892
rect 31556 73836 31948 73892
rect 38434 73836 38444 73892
rect 38500 73836 39004 73892
rect 39060 73836 39676 73892
rect 39732 73836 39742 73892
rect 40562 73836 40572 73892
rect 40628 73836 41468 73892
rect 41524 73836 41534 73892
rect 43586 73836 43596 73892
rect 43652 73836 43820 73892
rect 43876 73836 43886 73892
rect 44146 73836 44156 73892
rect 44212 73836 46284 73892
rect 46340 73836 46350 73892
rect 48626 73836 48636 73892
rect 48692 73836 49980 73892
rect 50036 73836 51772 73892
rect 51828 73836 51838 73892
rect 54450 73836 54460 73892
rect 54516 73836 54908 73892
rect 54964 73836 54974 73892
rect 55318 73836 55356 73892
rect 55412 73836 55422 73892
rect 57138 73836 57148 73892
rect 57204 73836 60508 73892
rect 60564 73836 60574 73892
rect 31892 73780 31948 73836
rect 31892 73724 34188 73780
rect 34244 73724 42700 73780
rect 42756 73724 42766 73780
rect 42914 73724 42924 73780
rect 42980 73724 44268 73780
rect 44324 73724 44334 73780
rect 44706 73724 44716 73780
rect 44772 73724 44940 73780
rect 44996 73724 45948 73780
rect 46004 73724 50428 73780
rect 51212 73724 57484 73780
rect 57540 73724 57550 73780
rect 58594 73724 58604 73780
rect 58660 73724 60956 73780
rect 61012 73724 61022 73780
rect 19826 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20110 73724
rect 37538 73612 37548 73668
rect 37604 73612 37772 73668
rect 37828 73612 38780 73668
rect 38836 73612 38846 73668
rect 43362 73612 43372 73668
rect 43428 73612 46620 73668
rect 46676 73612 46686 73668
rect 50372 73556 50428 73724
rect 50546 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50830 73724
rect 36866 73500 36876 73556
rect 36932 73500 38892 73556
rect 38948 73500 38958 73556
rect 41010 73500 41020 73556
rect 41076 73500 44044 73556
rect 44100 73500 44110 73556
rect 45714 73500 45724 73556
rect 45780 73500 46172 73556
rect 46228 73500 47852 73556
rect 47908 73500 47918 73556
rect 50372 73500 50988 73556
rect 51044 73500 51054 73556
rect 51212 73444 51268 73724
rect 51538 73612 51548 73668
rect 51604 73612 52332 73668
rect 52388 73612 52398 73668
rect 55234 73612 55244 73668
rect 55300 73612 59836 73668
rect 59892 73612 59902 73668
rect 54114 73500 54124 73556
rect 54180 73500 55356 73556
rect 55412 73500 55422 73556
rect 56018 73500 56028 73556
rect 56084 73500 57820 73556
rect 57876 73500 57886 73556
rect 37874 73388 37884 73444
rect 37940 73388 38668 73444
rect 43474 73388 43484 73444
rect 43540 73388 44212 73444
rect 44594 73388 44604 73444
rect 44660 73388 45612 73444
rect 45668 73388 47180 73444
rect 47236 73388 47246 73444
rect 48850 73388 48860 73444
rect 48916 73388 49420 73444
rect 49476 73388 51268 73444
rect 51986 73388 51996 73444
rect 52052 73388 53116 73444
rect 53172 73388 53182 73444
rect 54898 73388 54908 73444
rect 54964 73388 55916 73444
rect 55972 73388 55982 73444
rect 38612 73332 38668 73388
rect 44156 73332 44212 73388
rect 37650 73276 37660 73332
rect 37716 73276 38444 73332
rect 38500 73276 38510 73332
rect 38612 73276 38892 73332
rect 38948 73276 40012 73332
rect 40068 73276 40078 73332
rect 40786 73276 40796 73332
rect 40852 73276 43148 73332
rect 43204 73276 43932 73332
rect 43988 73276 43998 73332
rect 44156 73276 46060 73332
rect 46116 73276 46126 73332
rect 46274 73276 46284 73332
rect 46340 73276 47068 73332
rect 47124 73276 49644 73332
rect 49700 73276 49710 73332
rect 50306 73276 50316 73332
rect 50372 73276 50428 73388
rect 56914 73276 56924 73332
rect 56980 73276 57708 73332
rect 57764 73276 57774 73332
rect 59266 73276 59276 73332
rect 59332 73276 60172 73332
rect 60228 73276 66892 73332
rect 66948 73276 66958 73332
rect 40562 73164 40572 73220
rect 40628 73164 42700 73220
rect 42756 73164 47180 73220
rect 47236 73164 47246 73220
rect 49410 73164 49420 73220
rect 49476 73164 50764 73220
rect 50820 73164 50830 73220
rect 55682 73164 55692 73220
rect 55748 73164 56252 73220
rect 56308 73164 56812 73220
rect 56868 73164 56878 73220
rect 35522 73052 35532 73108
rect 35588 73052 38668 73108
rect 41010 73052 41020 73108
rect 41076 73052 42924 73108
rect 42980 73052 42990 73108
rect 44930 73052 44940 73108
rect 44996 73052 46284 73108
rect 46340 73052 46844 73108
rect 46900 73052 46910 73108
rect 38612 72996 38668 73052
rect 36978 72940 36988 72996
rect 37044 72940 37548 72996
rect 37604 72940 37614 72996
rect 38612 72940 43372 72996
rect 43428 72940 43438 72996
rect 4466 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4750 72940
rect 35186 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35470 72940
rect 49868 72884 49924 73164
rect 51062 73052 51100 73108
rect 51156 73052 51166 73108
rect 56578 73052 56588 73108
rect 56644 73052 59276 73108
rect 59332 73052 59342 73108
rect 65906 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66190 72940
rect 38658 72828 38668 72884
rect 38724 72828 40012 72884
rect 40068 72828 40078 72884
rect 49858 72828 49868 72884
rect 49924 72828 49934 72884
rect 41010 72716 41020 72772
rect 41076 72716 44156 72772
rect 44212 72716 44222 72772
rect 50866 72716 50876 72772
rect 50932 72716 51772 72772
rect 51828 72716 51838 72772
rect 53554 72716 53564 72772
rect 53620 72716 54460 72772
rect 54516 72716 54908 72772
rect 54964 72716 54974 72772
rect 30370 72604 30380 72660
rect 30436 72604 31276 72660
rect 31332 72604 31836 72660
rect 31892 72604 31948 72660
rect 32004 72604 32014 72660
rect 34178 72604 34188 72660
rect 34244 72604 35420 72660
rect 35476 72604 35486 72660
rect 37426 72604 37436 72660
rect 37492 72604 40572 72660
rect 40628 72604 41132 72660
rect 41188 72604 41692 72660
rect 41748 72604 41758 72660
rect 43138 72604 43148 72660
rect 43204 72604 45500 72660
rect 45556 72604 45566 72660
rect 49634 72604 49644 72660
rect 49700 72604 51548 72660
rect 51604 72604 51614 72660
rect 51986 72604 51996 72660
rect 52052 72604 53340 72660
rect 53396 72604 57148 72660
rect 57204 72604 57214 72660
rect 57474 72604 57484 72660
rect 57540 72604 59724 72660
rect 59780 72604 59790 72660
rect 37874 72492 37884 72548
rect 37940 72492 38444 72548
rect 38500 72492 40348 72548
rect 40404 72492 40414 72548
rect 41458 72492 41468 72548
rect 41524 72492 45164 72548
rect 45220 72492 46452 72548
rect 46610 72492 46620 72548
rect 46676 72492 47292 72548
rect 47348 72492 47358 72548
rect 47730 72492 47740 72548
rect 47796 72492 48412 72548
rect 48468 72492 48478 72548
rect 50082 72492 50092 72548
rect 50148 72492 50764 72548
rect 50820 72492 50830 72548
rect 51874 72492 51884 72548
rect 51940 72492 51950 72548
rect 52098 72492 52108 72548
rect 52164 72492 52444 72548
rect 52500 72492 53004 72548
rect 53060 72492 53070 72548
rect 53218 72492 53228 72548
rect 53284 72492 54684 72548
rect 54740 72492 58828 72548
rect 58884 72492 58894 72548
rect 46396 72436 46452 72492
rect 47740 72436 47796 72492
rect 36418 72380 36428 72436
rect 36484 72380 39228 72436
rect 39284 72380 39294 72436
rect 43586 72380 43596 72436
rect 43652 72380 43932 72436
rect 43988 72380 45052 72436
rect 45108 72380 45118 72436
rect 46386 72380 46396 72436
rect 46452 72380 47796 72436
rect 51884 72324 51940 72492
rect 52658 72380 52668 72436
rect 52724 72380 54348 72436
rect 54404 72380 54414 72436
rect 57026 72380 57036 72436
rect 57092 72380 59164 72436
rect 59220 72380 59230 72436
rect 15810 72268 15820 72324
rect 15876 72268 35308 72324
rect 35364 72268 35374 72324
rect 38546 72268 38556 72324
rect 38612 72268 39004 72324
rect 39060 72268 40012 72324
rect 40068 72268 41692 72324
rect 41748 72268 44604 72324
rect 44660 72268 44670 72324
rect 46274 72268 46284 72324
rect 46340 72268 47628 72324
rect 47684 72268 47694 72324
rect 49858 72268 49868 72324
rect 49924 72268 50316 72324
rect 50372 72268 50382 72324
rect 50978 72268 50988 72324
rect 51044 72268 51548 72324
rect 51604 72268 52892 72324
rect 52948 72268 54124 72324
rect 54180 72268 54190 72324
rect 19826 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20110 72156
rect 50546 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50830 72156
rect 56690 72044 56700 72100
rect 56756 72044 58716 72100
rect 58772 72044 60396 72100
rect 60452 72044 60462 72100
rect 36418 71932 36428 71988
rect 36484 71932 37772 71988
rect 37828 71932 37838 71988
rect 38770 71932 38780 71988
rect 38836 71932 39228 71988
rect 39284 71932 39294 71988
rect 46498 71932 46508 71988
rect 46564 71932 47852 71988
rect 47908 71932 48076 71988
rect 48132 71932 48142 71988
rect 59266 71932 59276 71988
rect 59332 71932 61404 71988
rect 61460 71932 61470 71988
rect 40114 71820 40124 71876
rect 40180 71820 41020 71876
rect 41076 71820 41086 71876
rect 42914 71820 42924 71876
rect 42980 71820 43260 71876
rect 43316 71820 45164 71876
rect 45220 71820 45230 71876
rect 55234 71820 55244 71876
rect 55300 71820 56700 71876
rect 56756 71820 56766 71876
rect 57362 71820 57372 71876
rect 57428 71820 57932 71876
rect 57988 71820 58940 71876
rect 58996 71820 59006 71876
rect 38770 71708 38780 71764
rect 38836 71708 39004 71764
rect 39060 71708 39070 71764
rect 41794 71708 41804 71764
rect 41860 71708 44492 71764
rect 44548 71708 44558 71764
rect 50194 71708 50204 71764
rect 50260 71708 51884 71764
rect 51940 71708 51950 71764
rect 41122 71596 41132 71652
rect 41188 71596 42252 71652
rect 42308 71596 42812 71652
rect 42868 71596 42878 71652
rect 42812 71540 42868 71596
rect 13794 71484 13804 71540
rect 13860 71484 34860 71540
rect 34916 71484 34926 71540
rect 38994 71484 39004 71540
rect 39060 71484 40124 71540
rect 40180 71484 40190 71540
rect 42812 71484 44940 71540
rect 44996 71484 45006 71540
rect 43586 71372 43596 71428
rect 43652 71372 44716 71428
rect 44772 71372 44782 71428
rect 4466 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4750 71372
rect 35186 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35470 71372
rect 65906 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66190 71372
rect 36194 71260 36204 71316
rect 36260 71260 48412 71316
rect 48468 71260 48478 71316
rect 39890 71148 39900 71204
rect 39956 71148 40348 71204
rect 40404 71148 41244 71204
rect 41300 71148 41310 71204
rect 46050 71148 46060 71204
rect 46116 71148 46396 71204
rect 46452 71148 46462 71204
rect 56130 71148 56140 71204
rect 56196 71148 57372 71204
rect 57428 71148 57438 71204
rect 34290 71036 34300 71092
rect 34356 71036 35196 71092
rect 35252 71036 35644 71092
rect 35700 71036 35710 71092
rect 38210 71036 38220 71092
rect 38276 71036 39004 71092
rect 39060 71036 39070 71092
rect 40226 71036 40236 71092
rect 40292 71036 40908 71092
rect 40964 71036 41804 71092
rect 41860 71036 41870 71092
rect 45042 71036 45052 71092
rect 45108 71036 45612 71092
rect 45668 71036 45678 71092
rect 47842 71036 47852 71092
rect 47908 71036 48748 71092
rect 48804 71036 48814 71092
rect 49298 71036 49308 71092
rect 49364 71036 50876 71092
rect 50932 71036 50942 71092
rect 51100 71036 73052 71092
rect 73108 71036 73118 71092
rect 48748 70980 48804 71036
rect 51100 70980 51156 71036
rect 36082 70924 36092 70980
rect 36148 70924 36428 70980
rect 36484 70924 38108 70980
rect 38164 70924 38174 70980
rect 39218 70924 39228 70980
rect 39284 70924 42812 70980
rect 42868 70924 42878 70980
rect 44818 70924 44828 70980
rect 44884 70924 46172 70980
rect 46228 70924 46238 70980
rect 48748 70924 51156 70980
rect 55458 70924 55468 70980
rect 55524 70924 55916 70980
rect 55972 70924 57036 70980
rect 57092 70924 57102 70980
rect 37762 70812 37772 70868
rect 37828 70812 39676 70868
rect 39732 70812 39742 70868
rect 39890 70700 39900 70756
rect 39956 70700 41020 70756
rect 41076 70700 41086 70756
rect 55234 70700 55244 70756
rect 55300 70700 55468 70756
rect 55524 70700 55534 70756
rect 38994 70588 39004 70644
rect 39060 70588 39788 70644
rect 39844 70588 39854 70644
rect 19826 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20110 70588
rect 50546 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50830 70588
rect 35522 70476 35532 70532
rect 35588 70476 45276 70532
rect 45332 70476 45342 70532
rect 52546 70476 52556 70532
rect 52612 70476 54572 70532
rect 54628 70476 55356 70532
rect 55412 70476 55422 70532
rect 31826 70364 31836 70420
rect 31892 70308 31948 70420
rect 36754 70364 36764 70420
rect 36820 70364 40124 70420
rect 40180 70364 40190 70420
rect 46162 70364 46172 70420
rect 46228 70364 48300 70420
rect 48356 70364 48366 70420
rect 50194 70364 50204 70420
rect 50260 70364 50652 70420
rect 50708 70364 50718 70420
rect 51650 70364 51660 70420
rect 51716 70364 53004 70420
rect 53060 70364 53070 70420
rect 54226 70364 54236 70420
rect 54292 70364 55468 70420
rect 55570 70364 55580 70420
rect 55636 70364 56028 70420
rect 56084 70364 56476 70420
rect 56532 70364 56542 70420
rect 55412 70308 55468 70364
rect 31892 70252 54124 70308
rect 54180 70252 54190 70308
rect 55412 70252 56588 70308
rect 56644 70252 56924 70308
rect 56980 70252 56990 70308
rect 36530 70140 36540 70196
rect 36596 70140 37212 70196
rect 37268 70140 37278 70196
rect 37538 70140 37548 70196
rect 37604 70140 39228 70196
rect 39284 70140 40124 70196
rect 40180 70140 40190 70196
rect 53442 70028 53452 70084
rect 53508 70028 55580 70084
rect 55636 70028 55646 70084
rect 4466 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4750 69804
rect 35186 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35470 69804
rect 65906 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66190 69804
rect 19826 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20110 69020
rect 50546 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50830 69020
rect 4466 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4750 68236
rect 35186 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35470 68236
rect 65906 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66190 68236
rect 19826 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20110 67452
rect 50546 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50830 67452
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 35186 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35470 66668
rect 65906 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66190 66668
rect 19826 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20110 65884
rect 50546 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50830 65884
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 35186 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35470 65100
rect 65906 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66190 65100
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 50546 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50830 64316
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 65906 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66190 63532
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 50546 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50830 62748
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 65906 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66190 61964
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 50546 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50830 61180
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 65906 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66190 60396
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 50546 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50830 59612
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 65906 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66190 58828
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 50546 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50830 58044
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 65906 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66190 57260
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 65906 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66190 55692
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 65906 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66190 54124
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 65906 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66190 52556
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 65906 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66190 50988
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 65906 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66190 49420
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 65906 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66190 47852
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 65906 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66190 46284
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 65906 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66190 44716
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 65906 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66190 43148
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 65906 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66190 41580
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 65906 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66190 40012
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 65906 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66190 38444
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 65906 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66190 36876
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 65906 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66190 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 65906 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66190 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 65906 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66190 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 65906 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66190 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 65906 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66190 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 65906 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66190 27468
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 65906 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66190 25900
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 65906 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66190 24332
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 65906 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66190 22764
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 65906 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66190 21196
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 65906 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66190 19628
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 65906 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66190 18060
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 65906 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66190 16492
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 65906 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66190 14924
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 65906 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66190 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 65906 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66190 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 65906 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66190 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 65906 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66190 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 65906 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66190 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 65906 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66190 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 65906 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66190 3948
rect 41794 3276 41804 3332
rect 41860 3276 42364 3332
rect 42420 3276 42430 3332
rect 43138 3276 43148 3332
rect 43204 3276 43708 3332
rect 43764 3276 43774 3332
rect 45154 3276 45164 3332
rect 45220 3276 45724 3332
rect 45780 3276 45790 3332
rect 46498 3276 46508 3332
rect 46564 3276 47068 3332
rect 47124 3276 47134 3332
rect 48514 3276 48524 3332
rect 48580 3276 49084 3332
rect 49140 3276 49150 3332
rect 49858 3276 49868 3332
rect 49924 3276 50428 3332
rect 50484 3276 50494 3332
rect 51874 3276 51884 3332
rect 51940 3276 52444 3332
rect 52500 3276 52510 3332
rect 53218 3276 53228 3332
rect 53284 3276 53788 3332
rect 53844 3276 53854 3332
rect 56578 3276 56588 3332
rect 56644 3276 57148 3332
rect 57204 3276 57214 3332
rect 58594 3276 58604 3332
rect 58660 3276 59164 3332
rect 59220 3276 59230 3332
rect 59938 3276 59948 3332
rect 60004 3276 60508 3332
rect 60564 3276 60574 3332
rect 61170 3276 61180 3332
rect 61236 3276 62300 3332
rect 62356 3276 62366 3332
rect 63186 3276 63196 3332
rect 63252 3276 64316 3332
rect 64372 3276 64382 3332
rect 64530 3276 64540 3332
rect 64596 3276 65660 3332
rect 65716 3276 65726 3332
rect 66546 3276 66556 3332
rect 66612 3276 67676 3332
rect 67732 3276 67742 3332
rect 67890 3276 67900 3332
rect 67956 3276 69020 3332
rect 69076 3276 69086 3332
rect 69906 3276 69916 3332
rect 69972 3276 71036 3332
rect 71092 3276 71102 3332
rect 71250 3276 71260 3332
rect 71316 3276 72380 3332
rect 72436 3276 72446 3332
rect 73378 3276 73388 3332
rect 73444 3276 74396 3332
rect 74452 3276 74462 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 55122 1708 55132 1764
rect 55188 1708 55804 1764
rect 55860 1708 55870 1764
rect 61842 1708 61852 1764
rect 61908 1708 62972 1764
rect 63028 1708 63038 1764
rect 65202 1708 65212 1764
rect 65268 1708 66332 1764
rect 66388 1708 66398 1764
rect 68562 1708 68572 1764
rect 68628 1708 69692 1764
rect 69748 1708 69758 1764
rect 71922 1708 71932 1764
rect 71988 1708 73052 1764
rect 73108 1708 73118 1764
<< via3 >>
rect 19836 76804 19892 76860
rect 19940 76804 19996 76860
rect 20044 76804 20100 76860
rect 50556 76804 50612 76860
rect 50660 76804 50716 76860
rect 50764 76804 50820 76860
rect 60284 76300 60340 76356
rect 60172 76076 60228 76132
rect 4476 76020 4532 76076
rect 4580 76020 4636 76076
rect 4684 76020 4740 76076
rect 35196 76020 35252 76076
rect 35300 76020 35356 76076
rect 35404 76020 35460 76076
rect 65916 76020 65972 76076
rect 66020 76020 66076 76076
rect 66124 76020 66180 76076
rect 39900 75740 39956 75796
rect 51100 75740 51156 75796
rect 55356 75628 55412 75684
rect 39900 75516 39956 75572
rect 32284 75404 32340 75460
rect 38612 75404 38668 75460
rect 43708 75404 43764 75460
rect 19836 75236 19892 75292
rect 19940 75236 19996 75292
rect 20044 75236 20100 75292
rect 50556 75236 50612 75292
rect 50660 75236 50716 75292
rect 50764 75236 50820 75292
rect 38668 75068 38724 75124
rect 55244 75068 55300 75124
rect 49756 74956 49812 75012
rect 43708 74844 43764 74900
rect 32284 74732 32340 74788
rect 49756 74732 49812 74788
rect 51548 74732 51604 74788
rect 4476 74452 4532 74508
rect 4580 74452 4636 74508
rect 4684 74452 4740 74508
rect 35196 74452 35252 74508
rect 35300 74452 35356 74508
rect 35404 74452 35460 74508
rect 65916 74452 65972 74508
rect 66020 74452 66076 74508
rect 66124 74452 66180 74508
rect 43484 74284 43540 74340
rect 43596 74172 43652 74228
rect 50988 74060 51044 74116
rect 51548 74060 51604 74116
rect 44604 73948 44660 74004
rect 51100 73948 51156 74004
rect 43596 73836 43652 73892
rect 55356 73836 55412 73892
rect 19836 73668 19892 73724
rect 19940 73668 19996 73724
rect 20044 73668 20100 73724
rect 50556 73668 50612 73724
rect 50660 73668 50716 73724
rect 50764 73668 50820 73724
rect 50988 73500 51044 73556
rect 55244 73612 55300 73668
rect 43484 73388 43540 73444
rect 4476 72884 4532 72940
rect 4580 72884 4636 72940
rect 4684 72884 4740 72940
rect 35196 72884 35252 72940
rect 35300 72884 35356 72940
rect 35404 72884 35460 72940
rect 51100 73052 51156 73108
rect 65916 72884 65972 72940
rect 66020 72884 66076 72940
rect 66124 72884 66180 72940
rect 44604 72268 44660 72324
rect 19836 72100 19892 72156
rect 19940 72100 19996 72156
rect 20044 72100 20100 72156
rect 50556 72100 50612 72156
rect 50660 72100 50716 72156
rect 50764 72100 50820 72156
rect 4476 71316 4532 71372
rect 4580 71316 4636 71372
rect 4684 71316 4740 71372
rect 35196 71316 35252 71372
rect 35300 71316 35356 71372
rect 35404 71316 35460 71372
rect 65916 71316 65972 71372
rect 66020 71316 66076 71372
rect 66124 71316 66180 71372
rect 19836 70532 19892 70588
rect 19940 70532 19996 70588
rect 20044 70532 20100 70588
rect 50556 70532 50612 70588
rect 50660 70532 50716 70588
rect 50764 70532 50820 70588
rect 4476 69748 4532 69804
rect 4580 69748 4636 69804
rect 4684 69748 4740 69804
rect 35196 69748 35252 69804
rect 35300 69748 35356 69804
rect 35404 69748 35460 69804
rect 65916 69748 65972 69804
rect 66020 69748 66076 69804
rect 66124 69748 66180 69804
rect 19836 68964 19892 69020
rect 19940 68964 19996 69020
rect 20044 68964 20100 69020
rect 50556 68964 50612 69020
rect 50660 68964 50716 69020
rect 50764 68964 50820 69020
rect 4476 68180 4532 68236
rect 4580 68180 4636 68236
rect 4684 68180 4740 68236
rect 35196 68180 35252 68236
rect 35300 68180 35356 68236
rect 35404 68180 35460 68236
rect 65916 68180 65972 68236
rect 66020 68180 66076 68236
rect 66124 68180 66180 68236
rect 19836 67396 19892 67452
rect 19940 67396 19996 67452
rect 20044 67396 20100 67452
rect 50556 67396 50612 67452
rect 50660 67396 50716 67452
rect 50764 67396 50820 67452
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 35196 66612 35252 66668
rect 35300 66612 35356 66668
rect 35404 66612 35460 66668
rect 65916 66612 65972 66668
rect 66020 66612 66076 66668
rect 66124 66612 66180 66668
rect 19836 65828 19892 65884
rect 19940 65828 19996 65884
rect 20044 65828 20100 65884
rect 50556 65828 50612 65884
rect 50660 65828 50716 65884
rect 50764 65828 50820 65884
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 35196 65044 35252 65100
rect 35300 65044 35356 65100
rect 35404 65044 35460 65100
rect 65916 65044 65972 65100
rect 66020 65044 66076 65100
rect 66124 65044 66180 65100
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 50556 64260 50612 64316
rect 50660 64260 50716 64316
rect 50764 64260 50820 64316
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 65916 63476 65972 63532
rect 66020 63476 66076 63532
rect 66124 63476 66180 63532
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 50556 62692 50612 62748
rect 50660 62692 50716 62748
rect 50764 62692 50820 62748
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 65916 61908 65972 61964
rect 66020 61908 66076 61964
rect 66124 61908 66180 61964
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 50556 61124 50612 61180
rect 50660 61124 50716 61180
rect 50764 61124 50820 61180
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 65916 60340 65972 60396
rect 66020 60340 66076 60396
rect 66124 60340 66180 60396
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 50556 59556 50612 59612
rect 50660 59556 50716 59612
rect 50764 59556 50820 59612
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 65916 58772 65972 58828
rect 66020 58772 66076 58828
rect 66124 58772 66180 58828
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 50556 57988 50612 58044
rect 50660 57988 50716 58044
rect 50764 57988 50820 58044
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 65916 57204 65972 57260
rect 66020 57204 66076 57260
rect 66124 57204 66180 57260
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 65916 55636 65972 55692
rect 66020 55636 66076 55692
rect 66124 55636 66180 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 65916 54068 65972 54124
rect 66020 54068 66076 54124
rect 66124 54068 66180 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 65916 52500 65972 52556
rect 66020 52500 66076 52556
rect 66124 52500 66180 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 65916 50932 65972 50988
rect 66020 50932 66076 50988
rect 66124 50932 66180 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 65916 49364 65972 49420
rect 66020 49364 66076 49420
rect 66124 49364 66180 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 65916 47796 65972 47852
rect 66020 47796 66076 47852
rect 66124 47796 66180 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 65916 46228 65972 46284
rect 66020 46228 66076 46284
rect 66124 46228 66180 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 65916 44660 65972 44716
rect 66020 44660 66076 44716
rect 66124 44660 66180 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 65916 43092 65972 43148
rect 66020 43092 66076 43148
rect 66124 43092 66180 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 65916 41524 65972 41580
rect 66020 41524 66076 41580
rect 66124 41524 66180 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 65916 39956 65972 40012
rect 66020 39956 66076 40012
rect 66124 39956 66180 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 65916 38388 65972 38444
rect 66020 38388 66076 38444
rect 66124 38388 66180 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 65916 36820 65972 36876
rect 66020 36820 66076 36876
rect 66124 36820 66180 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 65916 35252 65972 35308
rect 66020 35252 66076 35308
rect 66124 35252 66180 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 65916 33684 65972 33740
rect 66020 33684 66076 33740
rect 66124 33684 66180 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 65916 32116 65972 32172
rect 66020 32116 66076 32172
rect 66124 32116 66180 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 65916 30548 65972 30604
rect 66020 30548 66076 30604
rect 66124 30548 66180 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 65916 28980 65972 29036
rect 66020 28980 66076 29036
rect 66124 28980 66180 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 65916 27412 65972 27468
rect 66020 27412 66076 27468
rect 66124 27412 66180 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 65916 25844 65972 25900
rect 66020 25844 66076 25900
rect 66124 25844 66180 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 65916 24276 65972 24332
rect 66020 24276 66076 24332
rect 66124 24276 66180 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 65916 22708 65972 22764
rect 66020 22708 66076 22764
rect 66124 22708 66180 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 65916 21140 65972 21196
rect 66020 21140 66076 21196
rect 66124 21140 66180 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 65916 19572 65972 19628
rect 66020 19572 66076 19628
rect 66124 19572 66180 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 65916 18004 65972 18060
rect 66020 18004 66076 18060
rect 66124 18004 66180 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 65916 16436 65972 16492
rect 66020 16436 66076 16492
rect 66124 16436 66180 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 65916 14868 65972 14924
rect 66020 14868 66076 14924
rect 66124 14868 66180 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 65916 13300 65972 13356
rect 66020 13300 66076 13356
rect 66124 13300 66180 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 65916 11732 65972 11788
rect 66020 11732 66076 11788
rect 66124 11732 66180 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 65916 10164 65972 10220
rect 66020 10164 66076 10220
rect 66124 10164 66180 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 65916 8596 65972 8652
rect 66020 8596 66076 8652
rect 66124 8596 66180 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 65916 7028 65972 7084
rect 66020 7028 66076 7084
rect 66124 7028 66180 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 65916 5460 65972 5516
rect 66020 5460 66076 5516
rect 66124 5460 66180 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 65916 3892 65972 3948
rect 66020 3892 66076 3948
rect 66124 3892 66180 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 76076 4768 76892
rect 4448 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4768 76076
rect 4448 74508 4768 76020
rect 4448 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4768 74508
rect 4448 72940 4768 74452
rect 4448 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4768 72940
rect 4448 71372 4768 72884
rect 4448 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4768 71372
rect 4448 69804 4768 71316
rect 4448 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4768 69804
rect 4448 68236 4768 69748
rect 4448 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4768 68236
rect 4448 66668 4768 68180
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 76860 20128 76892
rect 19808 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20128 76860
rect 19808 75292 20128 76804
rect 35168 76076 35488 76892
rect 35168 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35488 76076
rect 19808 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20128 75292
rect 19808 73724 20128 75236
rect 32284 75460 32340 75470
rect 32284 74788 32340 75404
rect 32284 74722 32340 74732
rect 19808 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20128 73724
rect 19808 72156 20128 73668
rect 19808 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20128 72156
rect 19808 70588 20128 72100
rect 19808 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20128 70588
rect 19808 69020 20128 70532
rect 19808 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20128 69020
rect 19808 67452 20128 68964
rect 19808 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20128 67452
rect 19808 65884 20128 67396
rect 19808 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20128 65884
rect 19808 64316 20128 65828
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 19808 61180 20128 62692
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19808 56476 20128 57988
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 74508 35488 76020
rect 50528 76860 50848 76892
rect 50528 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50848 76860
rect 39900 75796 39956 75806
rect 39900 75572 39956 75740
rect 39900 75506 39956 75516
rect 38612 75460 38668 75470
rect 43708 75460 43764 75470
rect 38668 75404 38724 75460
rect 38612 75394 38724 75404
rect 38668 75124 38724 75394
rect 38668 75058 38724 75068
rect 43708 74900 43764 75404
rect 50528 75292 50848 76804
rect 60284 76356 60340 76366
rect 60172 76300 60284 76356
rect 60172 76132 60228 76300
rect 60284 76290 60340 76300
rect 60172 76066 60228 76076
rect 65888 76076 66208 76892
rect 65888 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66208 76076
rect 50528 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50848 75292
rect 43708 74834 43764 74844
rect 49756 75012 49812 75022
rect 49756 74788 49812 74956
rect 49756 74722 49812 74732
rect 35168 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35488 74508
rect 35168 72940 35488 74452
rect 43484 74340 43540 74350
rect 43484 73444 43540 74284
rect 43596 74228 43652 74238
rect 43596 73892 43652 74172
rect 43596 73826 43652 73836
rect 44604 74004 44660 74014
rect 43484 73378 43540 73388
rect 35168 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35488 72940
rect 35168 71372 35488 72884
rect 44604 72324 44660 73948
rect 44604 72258 44660 72268
rect 50528 73724 50848 75236
rect 51100 75796 51156 75806
rect 50528 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50848 73724
rect 35168 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35488 71372
rect 35168 69804 35488 71316
rect 35168 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35488 69804
rect 35168 68236 35488 69748
rect 35168 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35488 68236
rect 35168 66668 35488 68180
rect 35168 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35488 66668
rect 35168 65100 35488 66612
rect 35168 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35488 65100
rect 35168 63532 35488 65044
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 35168 61964 35488 63476
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 35168 60396 35488 61908
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 35168 57260 35488 58772
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 72156 50848 73668
rect 50988 74116 51044 74126
rect 50988 73556 51044 74060
rect 50988 73490 51044 73500
rect 51100 74004 51156 75740
rect 55356 75684 55412 75694
rect 55244 75124 55300 75134
rect 51548 74788 51604 74798
rect 51548 74116 51604 74732
rect 51548 74050 51604 74060
rect 51100 73108 51156 73948
rect 55244 73668 55300 75068
rect 55356 73892 55412 75628
rect 55356 73826 55412 73836
rect 65888 74508 66208 76020
rect 65888 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66208 74508
rect 55244 73602 55300 73612
rect 51100 73042 51156 73052
rect 50528 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50848 72156
rect 50528 70588 50848 72100
rect 50528 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50848 70588
rect 50528 69020 50848 70532
rect 50528 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50848 69020
rect 50528 67452 50848 68964
rect 50528 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50848 67452
rect 50528 65884 50848 67396
rect 50528 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50848 65884
rect 50528 64316 50848 65828
rect 50528 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50848 64316
rect 50528 62748 50848 64260
rect 50528 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50848 62748
rect 50528 61180 50848 62692
rect 50528 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50848 61180
rect 50528 59612 50848 61124
rect 50528 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50848 59612
rect 50528 58044 50848 59556
rect 50528 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50848 58044
rect 50528 56476 50848 57988
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 65888 72940 66208 74452
rect 65888 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66208 72940
rect 65888 71372 66208 72884
rect 65888 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66208 71372
rect 65888 69804 66208 71316
rect 65888 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66208 69804
rect 65888 68236 66208 69748
rect 65888 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66208 68236
rect 65888 66668 66208 68180
rect 65888 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66208 66668
rect 65888 65100 66208 66612
rect 65888 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66208 65100
rect 65888 63532 66208 65044
rect 65888 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66208 63532
rect 65888 61964 66208 63476
rect 65888 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66208 61964
rect 65888 60396 66208 61908
rect 65888 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66208 60396
rect 65888 58828 66208 60340
rect 65888 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66208 58828
rect 65888 57260 66208 58772
rect 65888 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66208 57260
rect 65888 55692 66208 57204
rect 65888 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66208 55692
rect 65888 54124 66208 55636
rect 65888 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66208 54124
rect 65888 52556 66208 54068
rect 65888 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66208 52556
rect 65888 50988 66208 52500
rect 65888 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66208 50988
rect 65888 49420 66208 50932
rect 65888 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66208 49420
rect 65888 47852 66208 49364
rect 65888 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66208 47852
rect 65888 46284 66208 47796
rect 65888 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66208 46284
rect 65888 44716 66208 46228
rect 65888 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66208 44716
rect 65888 43148 66208 44660
rect 65888 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66208 43148
rect 65888 41580 66208 43092
rect 65888 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66208 41580
rect 65888 40012 66208 41524
rect 65888 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66208 40012
rect 65888 38444 66208 39956
rect 65888 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66208 38444
rect 65888 36876 66208 38388
rect 65888 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66208 36876
rect 65888 35308 66208 36820
rect 65888 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66208 35308
rect 65888 33740 66208 35252
rect 65888 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66208 33740
rect 65888 32172 66208 33684
rect 65888 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66208 32172
rect 65888 30604 66208 32116
rect 65888 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66208 30604
rect 65888 29036 66208 30548
rect 65888 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66208 29036
rect 65888 27468 66208 28980
rect 65888 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66208 27468
rect 65888 25900 66208 27412
rect 65888 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66208 25900
rect 65888 24332 66208 25844
rect 65888 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66208 24332
rect 65888 22764 66208 24276
rect 65888 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66208 22764
rect 65888 21196 66208 22708
rect 65888 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66208 21196
rect 65888 19628 66208 21140
rect 65888 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66208 19628
rect 65888 18060 66208 19572
rect 65888 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66208 18060
rect 65888 16492 66208 18004
rect 65888 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66208 16492
rect 65888 14924 66208 16436
rect 65888 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66208 14924
rect 65888 13356 66208 14868
rect 65888 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66208 13356
rect 65888 11788 66208 13300
rect 65888 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66208 11788
rect 65888 10220 66208 11732
rect 65888 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66208 10220
rect 65888 8652 66208 10164
rect 65888 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66208 8652
rect 65888 7084 66208 8596
rect 65888 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66208 7084
rect 65888 5516 66208 7028
rect 65888 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66208 5516
rect 65888 3948 66208 5460
rect 65888 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66208 3948
rect 65888 3076 66208 3892
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__119__I dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 48720 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__123__A1
timestamp 1669390400
transform 1 0 48272 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__124__A1
timestamp 1669390400
transform 1 0 46480 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__124__A2
timestamp 1669390400
transform 1 0 46704 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__124__A3
timestamp 1669390400
transform 1 0 47152 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__125__A1
timestamp 1669390400
transform 1 0 46032 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__126__A1
timestamp 1669390400
transform 1 0 47600 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__I
timestamp 1669390400
transform 1 0 48496 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__A2
timestamp 1669390400
transform 1 0 47376 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__B2
timestamp 1669390400
transform 1 0 47824 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__129__A1
timestamp 1669390400
transform 1 0 46928 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__I
timestamp 1669390400
transform -1 0 38304 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__133__A2
timestamp 1669390400
transform 1 0 48048 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__134__A2
timestamp 1669390400
transform -1 0 38640 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__135__A2
timestamp 1669390400
transform -1 0 38640 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__136__I
timestamp 1669390400
transform -1 0 38192 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__137__A2
timestamp 1669390400
transform 1 0 44240 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__138__A1
timestamp 1669390400
transform 1 0 40992 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__138__A3
timestamp 1669390400
transform 1 0 41664 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__139__B1
timestamp 1669390400
transform 1 0 41664 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__141__A1
timestamp 1669390400
transform 1 0 46256 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__142__A1
timestamp 1669390400
transform 1 0 47600 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__147__I
timestamp 1669390400
transform 1 0 62496 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__150__A1
timestamp 1669390400
transform 1 0 61824 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__152__A1
timestamp 1669390400
transform -1 0 57008 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__152__A2
timestamp 1669390400
transform -1 0 56560 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__152__A3
timestamp 1669390400
transform 1 0 61600 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__153__A1
timestamp 1669390400
transform -1 0 55440 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__154__A1
timestamp 1669390400
transform 1 0 58240 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__155__A1
timestamp 1669390400
transform 1 0 55328 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__156__I
timestamp 1669390400
transform 1 0 63840 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__157__A2
timestamp 1669390400
transform 1 0 60592 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__157__B2
timestamp 1669390400
transform 1 0 61376 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__158__A1
timestamp 1669390400
transform 1 0 60144 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__159__A1
timestamp 1669390400
transform 1 0 54432 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__161__I
timestamp 1669390400
transform -1 0 55552 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__162__A2
timestamp 1669390400
transform 1 0 62048 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__165__I
timestamp 1669390400
transform 1 0 63392 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__167__A1
timestamp 1669390400
transform 1 0 58688 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__A1
timestamp 1669390400
transform 1 0 54880 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__170__A1
timestamp 1669390400
transform -1 0 54208 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__171__A1
timestamp 1669390400
transform -1 0 53088 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__171__B
timestamp 1669390400
transform -1 0 52640 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__176__I
timestamp 1669390400
transform -1 0 31024 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__A2
timestamp 1669390400
transform -1 0 50960 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__A2
timestamp 1669390400
transform -1 0 46480 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__B1
timestamp 1669390400
transform -1 0 45360 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__B2
timestamp 1669390400
transform -1 0 43344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__I
timestamp 1669390400
transform 1 0 35392 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__I
timestamp 1669390400
transform -1 0 34272 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__A1
timestamp 1669390400
transform 1 0 36400 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__A2
timestamp 1669390400
transform -1 0 36064 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__A1
timestamp 1669390400
transform -1 0 45808 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__A2
timestamp 1669390400
transform -1 0 44576 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__I
timestamp 1669390400
transform -1 0 46256 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__A1
timestamp 1669390400
transform 1 0 44912 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__A1
timestamp 1669390400
transform -1 0 56112 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__A1
timestamp 1669390400
transform -1 0 53536 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__I
timestamp 1669390400
transform -1 0 58016 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__I
timestamp 1669390400
transform 1 0 29232 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__A2
timestamp 1669390400
transform 1 0 30352 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__A2
timestamp 1669390400
transform -1 0 32480 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__A1
timestamp 1669390400
transform -1 0 29904 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__A2
timestamp 1669390400
transform -1 0 32032 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__A1
timestamp 1669390400
transform -1 0 37408 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__A2
timestamp 1669390400
transform -1 0 39760 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__A2
timestamp 1669390400
transform 1 0 37632 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__I
timestamp 1669390400
transform -1 0 38640 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__I
timestamp 1669390400
transform -1 0 59360 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__S
timestamp 1669390400
transform 1 0 59696 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__A2
timestamp 1669390400
transform -1 0 32928 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__A1
timestamp 1669390400
transform -1 0 33376 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__A2
timestamp 1669390400
transform -1 0 32256 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__I
timestamp 1669390400
transform -1 0 36512 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__A1
timestamp 1669390400
transform -1 0 44016 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__C
timestamp 1669390400
transform -1 0 44912 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__A1
timestamp 1669390400
transform 1 0 47824 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__A2
timestamp 1669390400
transform -1 0 54768 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__C
timestamp 1669390400
transform -1 0 54320 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__A3
timestamp 1669390400
transform 1 0 54432 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__I
timestamp 1669390400
transform 1 0 33824 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__A2
timestamp 1669390400
transform -1 0 35728 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__A2
timestamp 1669390400
transform -1 0 35280 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__A1
timestamp 1669390400
transform 1 0 45584 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__A1
timestamp 1669390400
transform -1 0 41104 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__A2
timestamp 1669390400
transform -1 0 39088 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__A1
timestamp 1669390400
transform 1 0 41664 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__A2
timestamp 1669390400
transform 1 0 44800 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__B
timestamp 1669390400
transform -1 0 39984 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__I0
timestamp 1669390400
transform 1 0 37520 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__A1
timestamp 1669390400
transform -1 0 52976 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__A1
timestamp 1669390400
transform 1 0 53200 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__A1
timestamp 1669390400
transform -1 0 51744 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__B
timestamp 1669390400
transform -1 0 51408 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__S
timestamp 1669390400
transform 1 0 49616 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__A1
timestamp 1669390400
transform -1 0 50736 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__A1
timestamp 1669390400
transform -1 0 50288 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__C
timestamp 1669390400
transform -1 0 49392 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__245__A2
timestamp 1669390400
transform -1 0 40208 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__A2
timestamp 1669390400
transform -1 0 36176 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__B1
timestamp 1669390400
transform -1 0 37296 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__A2
timestamp 1669390400
transform -1 0 33824 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__I
timestamp 1669390400
transform -1 0 29008 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1669390400
transform -1 0 1904 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform -1 0 39088 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1669390400
transform 1 0 42112 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1669390400
transform 1 0 44800 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1669390400
transform -1 0 47264 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1669390400
transform -1 0 46704 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1669390400
transform -1 0 49840 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1669390400
transform -1 0 51184 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1669390400
transform 1 0 62384 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1669390400
transform -1 0 54768 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1669390400
transform 1 0 60928 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1669390400
transform 1 0 59584 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1669390400
transform 1 0 62944 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1669390400
transform -1 0 63616 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1669390400
transform -1 0 65296 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1669390400
transform -1 0 66864 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1669390400
transform 1 0 70448 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1669390400
transform -1 0 70896 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1669390400
transform -1 0 72912 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1669390400
transform 1 0 77392 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1669390400
transform 1 0 78064 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output22_I
timestamp 1669390400
transform -1 0 6608 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output24_I
timestamp 1669390400
transform 1 0 26768 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output31_I
timestamp 1669390400
transform 1 0 13776 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output32_I
timestamp 1669390400
transform 1 0 15792 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output33_I
timestamp 1669390400
transform 1 0 17808 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output34_I
timestamp 1669390400
transform 1 0 19824 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output35_I
timestamp 1669390400
transform 1 0 20944 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output36_I
timestamp 1669390400
transform -1 0 24080 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5152 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 6048 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 6496 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 6720 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53
timestamp 1669390400
transform 1 0 7280 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65
timestamp 1669390400
transform 1 0 8624 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73
timestamp 1669390400
transform 1 0 9520 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81
timestamp 1669390400
transform 1 0 10416 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87
timestamp 1669390400
transform 1 0 11088 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93
timestamp 1669390400
transform 1 0 11760 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_99
timestamp 1669390400
transform 1 0 12432 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_105
timestamp 1669390400
transform 1 0 13104 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_111
timestamp 1669390400
transform 1 0 13776 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_117
timestamp 1669390400
transform 1 0 14448 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_123
timestamp 1669390400
transform 1 0 15120 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_129
timestamp 1669390400
transform 1 0 15792 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_135
timestamp 1669390400
transform 1 0 16464 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_141
timestamp 1669390400
transform 1 0 17136 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_147
timestamp 1669390400
transform 1 0 17808 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_153
timestamp 1669390400
transform 1 0 18480 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_159
timestamp 1669390400
transform 1 0 19152 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_165
timestamp 1669390400
transform 1 0 19824 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_171
timestamp 1669390400
transform 1 0 20496 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_177
timestamp 1669390400
transform 1 0 21168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_180
timestamp 1669390400
transform 1 0 21504 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_185
timestamp 1669390400
transform 1 0 22064 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_191
timestamp 1669390400
transform 1 0 22736 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_197
timestamp 1669390400
transform 1 0 23408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_203
timestamp 1669390400
transform 1 0 24080 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_209
timestamp 1669390400
transform 1 0 24752 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_215
timestamp 1669390400
transform 1 0 25424 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_221
timestamp 1669390400
transform 1 0 26096 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_227
timestamp 1669390400
transform 1 0 26768 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_233
timestamp 1669390400
transform 1 0 27440 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_239
timestamp 1669390400
transform 1 0 28112 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_245
timestamp 1669390400
transform 1 0 28784 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_251
timestamp 1669390400
transform 1 0 29456 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_257
timestamp 1669390400
transform 1 0 30128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_263
timestamp 1669390400
transform 1 0 30800 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_269
timestamp 1669390400
transform 1 0 31472 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_275
timestamp 1669390400
transform 1 0 32144 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_281
timestamp 1669390400
transform 1 0 32816 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_287
timestamp 1669390400
transform 1 0 33488 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_293
timestamp 1669390400
transform 1 0 34160 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_299
timestamp 1669390400
transform 1 0 34832 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_305
timestamp 1669390400
transform 1 0 35504 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_311
timestamp 1669390400
transform 1 0 36176 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_317
timestamp 1669390400
transform 1 0 36848 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_323
timestamp 1669390400
transform 1 0 37520 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_329
timestamp 1669390400
transform 1 0 38192 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_335
timestamp 1669390400
transform 1 0 38864 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_341
timestamp 1669390400
transform 1 0 39536 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_347
timestamp 1669390400
transform 1 0 40208 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_353
timestamp 1669390400
transform 1 0 40880 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_355
timestamp 1669390400
transform 1 0 41104 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_358
timestamp 1669390400
transform 1 0 41440 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_363
timestamp 1669390400
transform 1 0 42000 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_369
timestamp 1669390400
transform 1 0 42672 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_375
timestamp 1669390400
transform 1 0 43344 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_381
timestamp 1669390400
transform 1 0 44016 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_387
timestamp 1669390400
transform 1 0 44688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_393
timestamp 1669390400
transform 1 0 45360 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_399
timestamp 1669390400
transform 1 0 46032 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_405
timestamp 1669390400
transform 1 0 46704 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_411
timestamp 1669390400
transform 1 0 47376 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_417
timestamp 1669390400
transform 1 0 48048 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_423
timestamp 1669390400
transform 1 0 48720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_429
timestamp 1669390400
transform 1 0 49392 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_435
timestamp 1669390400
transform 1 0 50064 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_441
timestamp 1669390400
transform 1 0 50736 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_447
timestamp 1669390400
transform 1 0 51408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_453
timestamp 1669390400
transform 1 0 52080 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_459
timestamp 1669390400
transform 1 0 52752 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_465
timestamp 1669390400
transform 1 0 53424 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_471
timestamp 1669390400
transform 1 0 54096 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_477
timestamp 1669390400
transform 1 0 54768 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_483
timestamp 1669390400
transform 1 0 55440 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_489
timestamp 1669390400
transform 1 0 56112 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_495
timestamp 1669390400
transform 1 0 56784 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_501
timestamp 1669390400
transform 1 0 57456 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_507
timestamp 1669390400
transform 1 0 58128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_513
timestamp 1669390400
transform 1 0 58800 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_519
timestamp 1669390400
transform 1 0 59472 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_525
timestamp 1669390400
transform 1 0 60144 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_531
timestamp 1669390400
transform 1 0 60816 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_533
timestamp 1669390400
transform 1 0 61040 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_536
timestamp 1669390400
transform 1 0 61376 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_541
timestamp 1669390400
transform 1 0 61936 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_547
timestamp 1669390400
transform 1 0 62608 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_553
timestamp 1669390400
transform 1 0 63280 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_559
timestamp 1669390400
transform 1 0 63952 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_565
timestamp 1669390400
transform 1 0 64624 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_571
timestamp 1669390400
transform 1 0 65296 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_577
timestamp 1669390400
transform 1 0 65968 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_583
timestamp 1669390400
transform 1 0 66640 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_589
timestamp 1669390400
transform 1 0 67312 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_595
timestamp 1669390400
transform 1 0 67984 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_601
timestamp 1669390400
transform 1 0 68656 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_607
timestamp 1669390400
transform 1 0 69328 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_613
timestamp 1669390400
transform 1 0 70000 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_619
timestamp 1669390400
transform 1 0 70672 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_625
timestamp 1669390400
transform 1 0 71344 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_631
timestamp 1669390400
transform 1 0 72016 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_637
timestamp 1669390400
transform 1 0 72688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_643
timestamp 1669390400
transform 1 0 73360 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_649
timestamp 1669390400
transform 1 0 74032 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_655
timestamp 1669390400
transform 1 0 74704 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_687
timestamp 1669390400
transform 1 0 78288 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_66
timestamp 1669390400
transform 1 0 8736 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_130
timestamp 1669390400
transform 1 0 15904 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_194
timestamp 1669390400
transform 1 0 23072 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_258
timestamp 1669390400
transform 1 0 30240 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_322
timestamp 1669390400
transform 1 0 37408 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_354
timestamp 1669390400
transform 1 0 40992 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_356
timestamp 1669390400
transform 1 0 41216 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_359
timestamp 1669390400
transform 1 0 41552 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_423
timestamp 1669390400
transform 1 0 48720 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_487
timestamp 1669390400
transform 1 0 55888 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_551
timestamp 1669390400
transform 1 0 63056 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_615 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 70224 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_631
timestamp 1669390400
transform 1 0 72016 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_639
timestamp 1669390400
transform 1 0 72912 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_645
timestamp 1669390400
transform 1 0 73584 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_651
timestamp 1669390400
transform 1 0 74256 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_683
timestamp 1669390400
transform 1 0 77840 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_687
timestamp 1669390400
transform 1 0 78288 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_2
timestamp 1669390400
transform 1 0 1568 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_66
timestamp 1669390400
transform 1 0 8736 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_130
timestamp 1669390400
transform 1 0 15904 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_162
timestamp 1669390400
transform 1 0 19488 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_180
timestamp 1669390400
transform 1 0 21504 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_244
timestamp 1669390400
transform 1 0 28672 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_308
timestamp 1669390400
transform 1 0 35840 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_372
timestamp 1669390400
transform 1 0 43008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_436
timestamp 1669390400
transform 1 0 50176 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_500
timestamp 1669390400
transform 1 0 57344 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_532
timestamp 1669390400
transform 1 0 60928 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_534
timestamp 1669390400
transform 1 0 61152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_537
timestamp 1669390400
transform 1 0 61488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_601
timestamp 1669390400
transform 1 0 68656 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_665
timestamp 1669390400
transform 1 0 75824 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_681
timestamp 1669390400
transform 1 0 77616 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_685
timestamp 1669390400
transform 1 0 78064 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_687
timestamp 1669390400
transform 1 0 78288 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1669390400
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_66
timestamp 1669390400
transform 1 0 8736 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_130
timestamp 1669390400
transform 1 0 15904 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_194
timestamp 1669390400
transform 1 0 23072 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_258
timestamp 1669390400
transform 1 0 30240 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_322
timestamp 1669390400
transform 1 0 37408 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_354
timestamp 1669390400
transform 1 0 40992 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_356
timestamp 1669390400
transform 1 0 41216 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_359
timestamp 1669390400
transform 1 0 41552 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_423
timestamp 1669390400
transform 1 0 48720 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_487
timestamp 1669390400
transform 1 0 55888 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_551
timestamp 1669390400
transform 1 0 63056 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_615
timestamp 1669390400
transform 1 0 70224 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_679
timestamp 1669390400
transform 1 0 77392 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_687
timestamp 1669390400
transform 1 0 78288 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_2
timestamp 1669390400
transform 1 0 1568 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_66
timestamp 1669390400
transform 1 0 8736 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_130
timestamp 1669390400
transform 1 0 15904 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_162
timestamp 1669390400
transform 1 0 19488 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_180
timestamp 1669390400
transform 1 0 21504 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_244
timestamp 1669390400
transform 1 0 28672 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_308
timestamp 1669390400
transform 1 0 35840 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_372
timestamp 1669390400
transform 1 0 43008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_436
timestamp 1669390400
transform 1 0 50176 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_500
timestamp 1669390400
transform 1 0 57344 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_532
timestamp 1669390400
transform 1 0 60928 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_534
timestamp 1669390400
transform 1 0 61152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_537
timestamp 1669390400
transform 1 0 61488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_601
timestamp 1669390400
transform 1 0 68656 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_665
timestamp 1669390400
transform 1 0 75824 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_681
timestamp 1669390400
transform 1 0 77616 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_685
timestamp 1669390400
transform 1 0 78064 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_687
timestamp 1669390400
transform 1 0 78288 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1669390400
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_66
timestamp 1669390400
transform 1 0 8736 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_130
timestamp 1669390400
transform 1 0 15904 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_194
timestamp 1669390400
transform 1 0 23072 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_258
timestamp 1669390400
transform 1 0 30240 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_322
timestamp 1669390400
transform 1 0 37408 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_354
timestamp 1669390400
transform 1 0 40992 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_356
timestamp 1669390400
transform 1 0 41216 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_359
timestamp 1669390400
transform 1 0 41552 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_423
timestamp 1669390400
transform 1 0 48720 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_487
timestamp 1669390400
transform 1 0 55888 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_551
timestamp 1669390400
transform 1 0 63056 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_615
timestamp 1669390400
transform 1 0 70224 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_679
timestamp 1669390400
transform 1 0 77392 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_687
timestamp 1669390400
transform 1 0 78288 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_2
timestamp 1669390400
transform 1 0 1568 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_66
timestamp 1669390400
transform 1 0 8736 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_130
timestamp 1669390400
transform 1 0 15904 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_162
timestamp 1669390400
transform 1 0 19488 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_180
timestamp 1669390400
transform 1 0 21504 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_244
timestamp 1669390400
transform 1 0 28672 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_308
timestamp 1669390400
transform 1 0 35840 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_372
timestamp 1669390400
transform 1 0 43008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_436
timestamp 1669390400
transform 1 0 50176 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_500
timestamp 1669390400
transform 1 0 57344 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_532
timestamp 1669390400
transform 1 0 60928 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_534
timestamp 1669390400
transform 1 0 61152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_537
timestamp 1669390400
transform 1 0 61488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_601
timestamp 1669390400
transform 1 0 68656 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_665
timestamp 1669390400
transform 1 0 75824 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_681
timestamp 1669390400
transform 1 0 77616 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_685
timestamp 1669390400
transform 1 0 78064 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_687
timestamp 1669390400
transform 1 0 78288 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1669390400
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_66
timestamp 1669390400
transform 1 0 8736 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_130
timestamp 1669390400
transform 1 0 15904 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_194
timestamp 1669390400
transform 1 0 23072 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_258
timestamp 1669390400
transform 1 0 30240 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_322
timestamp 1669390400
transform 1 0 37408 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_354
timestamp 1669390400
transform 1 0 40992 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_356
timestamp 1669390400
transform 1 0 41216 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_359
timestamp 1669390400
transform 1 0 41552 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_423
timestamp 1669390400
transform 1 0 48720 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_487
timestamp 1669390400
transform 1 0 55888 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_551
timestamp 1669390400
transform 1 0 63056 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_615
timestamp 1669390400
transform 1 0 70224 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_679
timestamp 1669390400
transform 1 0 77392 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_687
timestamp 1669390400
transform 1 0 78288 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_2
timestamp 1669390400
transform 1 0 1568 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_66
timestamp 1669390400
transform 1 0 8736 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_130
timestamp 1669390400
transform 1 0 15904 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_162
timestamp 1669390400
transform 1 0 19488 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_180
timestamp 1669390400
transform 1 0 21504 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_244
timestamp 1669390400
transform 1 0 28672 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_308
timestamp 1669390400
transform 1 0 35840 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_372
timestamp 1669390400
transform 1 0 43008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_436
timestamp 1669390400
transform 1 0 50176 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_500
timestamp 1669390400
transform 1 0 57344 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_532
timestamp 1669390400
transform 1 0 60928 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_534
timestamp 1669390400
transform 1 0 61152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_537
timestamp 1669390400
transform 1 0 61488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_601
timestamp 1669390400
transform 1 0 68656 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_665
timestamp 1669390400
transform 1 0 75824 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_681
timestamp 1669390400
transform 1 0 77616 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_685
timestamp 1669390400
transform 1 0 78064 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_687
timestamp 1669390400
transform 1 0 78288 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1669390400
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_66
timestamp 1669390400
transform 1 0 8736 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_130
timestamp 1669390400
transform 1 0 15904 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_194
timestamp 1669390400
transform 1 0 23072 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_258
timestamp 1669390400
transform 1 0 30240 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_322
timestamp 1669390400
transform 1 0 37408 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_354
timestamp 1669390400
transform 1 0 40992 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_356
timestamp 1669390400
transform 1 0 41216 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_359
timestamp 1669390400
transform 1 0 41552 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_423
timestamp 1669390400
transform 1 0 48720 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_487
timestamp 1669390400
transform 1 0 55888 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_551
timestamp 1669390400
transform 1 0 63056 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_615
timestamp 1669390400
transform 1 0 70224 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_679
timestamp 1669390400
transform 1 0 77392 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_687
timestamp 1669390400
transform 1 0 78288 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_2
timestamp 1669390400
transform 1 0 1568 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_66
timestamp 1669390400
transform 1 0 8736 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_130
timestamp 1669390400
transform 1 0 15904 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_162
timestamp 1669390400
transform 1 0 19488 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_180
timestamp 1669390400
transform 1 0 21504 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_244
timestamp 1669390400
transform 1 0 28672 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_308
timestamp 1669390400
transform 1 0 35840 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_372
timestamp 1669390400
transform 1 0 43008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_436
timestamp 1669390400
transform 1 0 50176 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_500
timestamp 1669390400
transform 1 0 57344 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_532
timestamp 1669390400
transform 1 0 60928 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_534
timestamp 1669390400
transform 1 0 61152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_537
timestamp 1669390400
transform 1 0 61488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_601
timestamp 1669390400
transform 1 0 68656 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_665
timestamp 1669390400
transform 1 0 75824 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_681
timestamp 1669390400
transform 1 0 77616 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_685
timestamp 1669390400
transform 1 0 78064 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_687
timestamp 1669390400
transform 1 0 78288 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1669390400
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_66
timestamp 1669390400
transform 1 0 8736 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_130
timestamp 1669390400
transform 1 0 15904 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_194
timestamp 1669390400
transform 1 0 23072 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_258
timestamp 1669390400
transform 1 0 30240 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_322
timestamp 1669390400
transform 1 0 37408 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_354
timestamp 1669390400
transform 1 0 40992 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_356
timestamp 1669390400
transform 1 0 41216 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_359
timestamp 1669390400
transform 1 0 41552 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_423
timestamp 1669390400
transform 1 0 48720 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_487
timestamp 1669390400
transform 1 0 55888 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_551
timestamp 1669390400
transform 1 0 63056 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_615
timestamp 1669390400
transform 1 0 70224 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_679
timestamp 1669390400
transform 1 0 77392 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_687
timestamp 1669390400
transform 1 0 78288 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_2
timestamp 1669390400
transform 1 0 1568 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_66
timestamp 1669390400
transform 1 0 8736 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_130
timestamp 1669390400
transform 1 0 15904 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_162
timestamp 1669390400
transform 1 0 19488 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_180
timestamp 1669390400
transform 1 0 21504 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_244
timestamp 1669390400
transform 1 0 28672 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_308
timestamp 1669390400
transform 1 0 35840 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_372
timestamp 1669390400
transform 1 0 43008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_436
timestamp 1669390400
transform 1 0 50176 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_500
timestamp 1669390400
transform 1 0 57344 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_532
timestamp 1669390400
transform 1 0 60928 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_534
timestamp 1669390400
transform 1 0 61152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_537
timestamp 1669390400
transform 1 0 61488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_601
timestamp 1669390400
transform 1 0 68656 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_665
timestamp 1669390400
transform 1 0 75824 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_681
timestamp 1669390400
transform 1 0 77616 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_685
timestamp 1669390400
transform 1 0 78064 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_687
timestamp 1669390400
transform 1 0 78288 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1669390400
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_66
timestamp 1669390400
transform 1 0 8736 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_130
timestamp 1669390400
transform 1 0 15904 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_194
timestamp 1669390400
transform 1 0 23072 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_258
timestamp 1669390400
transform 1 0 30240 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_322
timestamp 1669390400
transform 1 0 37408 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_354
timestamp 1669390400
transform 1 0 40992 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_356
timestamp 1669390400
transform 1 0 41216 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_359
timestamp 1669390400
transform 1 0 41552 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_423
timestamp 1669390400
transform 1 0 48720 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_487
timestamp 1669390400
transform 1 0 55888 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_551
timestamp 1669390400
transform 1 0 63056 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_615
timestamp 1669390400
transform 1 0 70224 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_679
timestamp 1669390400
transform 1 0 77392 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_687
timestamp 1669390400
transform 1 0 78288 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_2
timestamp 1669390400
transform 1 0 1568 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_66
timestamp 1669390400
transform 1 0 8736 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_130
timestamp 1669390400
transform 1 0 15904 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_162
timestamp 1669390400
transform 1 0 19488 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_180
timestamp 1669390400
transform 1 0 21504 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_244
timestamp 1669390400
transform 1 0 28672 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_308
timestamp 1669390400
transform 1 0 35840 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_372
timestamp 1669390400
transform 1 0 43008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_436
timestamp 1669390400
transform 1 0 50176 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_500
timestamp 1669390400
transform 1 0 57344 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_532
timestamp 1669390400
transform 1 0 60928 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_534
timestamp 1669390400
transform 1 0 61152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_537
timestamp 1669390400
transform 1 0 61488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_601
timestamp 1669390400
transform 1 0 68656 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_665
timestamp 1669390400
transform 1 0 75824 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_681
timestamp 1669390400
transform 1 0 77616 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_685
timestamp 1669390400
transform 1 0 78064 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_687
timestamp 1669390400
transform 1 0 78288 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1669390400
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_66
timestamp 1669390400
transform 1 0 8736 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_130
timestamp 1669390400
transform 1 0 15904 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_194
timestamp 1669390400
transform 1 0 23072 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_258
timestamp 1669390400
transform 1 0 30240 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_322
timestamp 1669390400
transform 1 0 37408 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_354
timestamp 1669390400
transform 1 0 40992 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_356
timestamp 1669390400
transform 1 0 41216 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_359
timestamp 1669390400
transform 1 0 41552 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_423
timestamp 1669390400
transform 1 0 48720 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_487
timestamp 1669390400
transform 1 0 55888 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_551
timestamp 1669390400
transform 1 0 63056 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_615
timestamp 1669390400
transform 1 0 70224 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_679
timestamp 1669390400
transform 1 0 77392 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_687
timestamp 1669390400
transform 1 0 78288 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_2
timestamp 1669390400
transform 1 0 1568 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_66
timestamp 1669390400
transform 1 0 8736 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_130
timestamp 1669390400
transform 1 0 15904 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_162
timestamp 1669390400
transform 1 0 19488 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_180
timestamp 1669390400
transform 1 0 21504 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_244
timestamp 1669390400
transform 1 0 28672 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_308
timestamp 1669390400
transform 1 0 35840 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_372
timestamp 1669390400
transform 1 0 43008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_436
timestamp 1669390400
transform 1 0 50176 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_500
timestamp 1669390400
transform 1 0 57344 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_532
timestamp 1669390400
transform 1 0 60928 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_534
timestamp 1669390400
transform 1 0 61152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_537
timestamp 1669390400
transform 1 0 61488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_601
timestamp 1669390400
transform 1 0 68656 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_665
timestamp 1669390400
transform 1 0 75824 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_681
timestamp 1669390400
transform 1 0 77616 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_685
timestamp 1669390400
transform 1 0 78064 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_687
timestamp 1669390400
transform 1 0 78288 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_2
timestamp 1669390400
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_66
timestamp 1669390400
transform 1 0 8736 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_130
timestamp 1669390400
transform 1 0 15904 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_194
timestamp 1669390400
transform 1 0 23072 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_258
timestamp 1669390400
transform 1 0 30240 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_322
timestamp 1669390400
transform 1 0 37408 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_354
timestamp 1669390400
transform 1 0 40992 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_356
timestamp 1669390400
transform 1 0 41216 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_359
timestamp 1669390400
transform 1 0 41552 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_423
timestamp 1669390400
transform 1 0 48720 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_487
timestamp 1669390400
transform 1 0 55888 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_551
timestamp 1669390400
transform 1 0 63056 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_615
timestamp 1669390400
transform 1 0 70224 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_679
timestamp 1669390400
transform 1 0 77392 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_687
timestamp 1669390400
transform 1 0 78288 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_2
timestamp 1669390400
transform 1 0 1568 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_66
timestamp 1669390400
transform 1 0 8736 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_130
timestamp 1669390400
transform 1 0 15904 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_162
timestamp 1669390400
transform 1 0 19488 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_180
timestamp 1669390400
transform 1 0 21504 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_244
timestamp 1669390400
transform 1 0 28672 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_308
timestamp 1669390400
transform 1 0 35840 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_372
timestamp 1669390400
transform 1 0 43008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_436
timestamp 1669390400
transform 1 0 50176 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_500
timestamp 1669390400
transform 1 0 57344 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_532
timestamp 1669390400
transform 1 0 60928 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_534
timestamp 1669390400
transform 1 0 61152 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_537
timestamp 1669390400
transform 1 0 61488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_601
timestamp 1669390400
transform 1 0 68656 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_665
timestamp 1669390400
transform 1 0 75824 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_681
timestamp 1669390400
transform 1 0 77616 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_685
timestamp 1669390400
transform 1 0 78064 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_687
timestamp 1669390400
transform 1 0 78288 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_2
timestamp 1669390400
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_66
timestamp 1669390400
transform 1 0 8736 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_130
timestamp 1669390400
transform 1 0 15904 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_194
timestamp 1669390400
transform 1 0 23072 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_258
timestamp 1669390400
transform 1 0 30240 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_322
timestamp 1669390400
transform 1 0 37408 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_354
timestamp 1669390400
transform 1 0 40992 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_356
timestamp 1669390400
transform 1 0 41216 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_359
timestamp 1669390400
transform 1 0 41552 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_423
timestamp 1669390400
transform 1 0 48720 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_487
timestamp 1669390400
transform 1 0 55888 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_551
timestamp 1669390400
transform 1 0 63056 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_615
timestamp 1669390400
transform 1 0 70224 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_679
timestamp 1669390400
transform 1 0 77392 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_687
timestamp 1669390400
transform 1 0 78288 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_2
timestamp 1669390400
transform 1 0 1568 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_66
timestamp 1669390400
transform 1 0 8736 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_130
timestamp 1669390400
transform 1 0 15904 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_162
timestamp 1669390400
transform 1 0 19488 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_180
timestamp 1669390400
transform 1 0 21504 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_244
timestamp 1669390400
transform 1 0 28672 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_308
timestamp 1669390400
transform 1 0 35840 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_372
timestamp 1669390400
transform 1 0 43008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_436
timestamp 1669390400
transform 1 0 50176 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_500
timestamp 1669390400
transform 1 0 57344 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_532
timestamp 1669390400
transform 1 0 60928 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_534
timestamp 1669390400
transform 1 0 61152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_537
timestamp 1669390400
transform 1 0 61488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_601
timestamp 1669390400
transform 1 0 68656 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_665
timestamp 1669390400
transform 1 0 75824 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_681
timestamp 1669390400
transform 1 0 77616 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_685
timestamp 1669390400
transform 1 0 78064 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_687
timestamp 1669390400
transform 1 0 78288 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1669390400
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_66
timestamp 1669390400
transform 1 0 8736 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_130
timestamp 1669390400
transform 1 0 15904 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_194
timestamp 1669390400
transform 1 0 23072 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_258
timestamp 1669390400
transform 1 0 30240 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_322
timestamp 1669390400
transform 1 0 37408 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_354
timestamp 1669390400
transform 1 0 40992 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_356
timestamp 1669390400
transform 1 0 41216 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_359
timestamp 1669390400
transform 1 0 41552 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_423
timestamp 1669390400
transform 1 0 48720 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_487
timestamp 1669390400
transform 1 0 55888 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_551
timestamp 1669390400
transform 1 0 63056 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_615
timestamp 1669390400
transform 1 0 70224 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_679
timestamp 1669390400
transform 1 0 77392 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_687
timestamp 1669390400
transform 1 0 78288 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_2
timestamp 1669390400
transform 1 0 1568 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_66
timestamp 1669390400
transform 1 0 8736 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_130
timestamp 1669390400
transform 1 0 15904 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_162
timestamp 1669390400
transform 1 0 19488 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_180
timestamp 1669390400
transform 1 0 21504 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_244
timestamp 1669390400
transform 1 0 28672 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_308
timestamp 1669390400
transform 1 0 35840 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_372
timestamp 1669390400
transform 1 0 43008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_436
timestamp 1669390400
transform 1 0 50176 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_500
timestamp 1669390400
transform 1 0 57344 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_532
timestamp 1669390400
transform 1 0 60928 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_534
timestamp 1669390400
transform 1 0 61152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_537
timestamp 1669390400
transform 1 0 61488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_601
timestamp 1669390400
transform 1 0 68656 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_665
timestamp 1669390400
transform 1 0 75824 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_681
timestamp 1669390400
transform 1 0 77616 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_685
timestamp 1669390400
transform 1 0 78064 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_687
timestamp 1669390400
transform 1 0 78288 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_2
timestamp 1669390400
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_66
timestamp 1669390400
transform 1 0 8736 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_130
timestamp 1669390400
transform 1 0 15904 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_194
timestamp 1669390400
transform 1 0 23072 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_258
timestamp 1669390400
transform 1 0 30240 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_322
timestamp 1669390400
transform 1 0 37408 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_354
timestamp 1669390400
transform 1 0 40992 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_356
timestamp 1669390400
transform 1 0 41216 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_359
timestamp 1669390400
transform 1 0 41552 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_423
timestamp 1669390400
transform 1 0 48720 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_487
timestamp 1669390400
transform 1 0 55888 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_551
timestamp 1669390400
transform 1 0 63056 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_615
timestamp 1669390400
transform 1 0 70224 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_679
timestamp 1669390400
transform 1 0 77392 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_687
timestamp 1669390400
transform 1 0 78288 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_2
timestamp 1669390400
transform 1 0 1568 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_66
timestamp 1669390400
transform 1 0 8736 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_130
timestamp 1669390400
transform 1 0 15904 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_162
timestamp 1669390400
transform 1 0 19488 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_180
timestamp 1669390400
transform 1 0 21504 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_244
timestamp 1669390400
transform 1 0 28672 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_308
timestamp 1669390400
transform 1 0 35840 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_372
timestamp 1669390400
transform 1 0 43008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_436
timestamp 1669390400
transform 1 0 50176 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_500
timestamp 1669390400
transform 1 0 57344 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_532
timestamp 1669390400
transform 1 0 60928 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_534
timestamp 1669390400
transform 1 0 61152 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_537
timestamp 1669390400
transform 1 0 61488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_601
timestamp 1669390400
transform 1 0 68656 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_665
timestamp 1669390400
transform 1 0 75824 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_681
timestamp 1669390400
transform 1 0 77616 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_685
timestamp 1669390400
transform 1 0 78064 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_687
timestamp 1669390400
transform 1 0 78288 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_2
timestamp 1669390400
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_66
timestamp 1669390400
transform 1 0 8736 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_130
timestamp 1669390400
transform 1 0 15904 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_194
timestamp 1669390400
transform 1 0 23072 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_258
timestamp 1669390400
transform 1 0 30240 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_322
timestamp 1669390400
transform 1 0 37408 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_354
timestamp 1669390400
transform 1 0 40992 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_356
timestamp 1669390400
transform 1 0 41216 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_359
timestamp 1669390400
transform 1 0 41552 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_423
timestamp 1669390400
transform 1 0 48720 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_487
timestamp 1669390400
transform 1 0 55888 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_551
timestamp 1669390400
transform 1 0 63056 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_615
timestamp 1669390400
transform 1 0 70224 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_679
timestamp 1669390400
transform 1 0 77392 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_687
timestamp 1669390400
transform 1 0 78288 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_2
timestamp 1669390400
transform 1 0 1568 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_66
timestamp 1669390400
transform 1 0 8736 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_130
timestamp 1669390400
transform 1 0 15904 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_162
timestamp 1669390400
transform 1 0 19488 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_180
timestamp 1669390400
transform 1 0 21504 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_244
timestamp 1669390400
transform 1 0 28672 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_308
timestamp 1669390400
transform 1 0 35840 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_372
timestamp 1669390400
transform 1 0 43008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_436
timestamp 1669390400
transform 1 0 50176 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_500
timestamp 1669390400
transform 1 0 57344 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_532
timestamp 1669390400
transform 1 0 60928 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_534
timestamp 1669390400
transform 1 0 61152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_537
timestamp 1669390400
transform 1 0 61488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_601
timestamp 1669390400
transform 1 0 68656 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_665
timestamp 1669390400
transform 1 0 75824 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_681
timestamp 1669390400
transform 1 0 77616 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_685
timestamp 1669390400
transform 1 0 78064 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_687
timestamp 1669390400
transform 1 0 78288 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_2
timestamp 1669390400
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_66
timestamp 1669390400
transform 1 0 8736 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_130
timestamp 1669390400
transform 1 0 15904 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_194
timestamp 1669390400
transform 1 0 23072 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_258
timestamp 1669390400
transform 1 0 30240 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_322
timestamp 1669390400
transform 1 0 37408 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_354
timestamp 1669390400
transform 1 0 40992 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_356
timestamp 1669390400
transform 1 0 41216 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_359
timestamp 1669390400
transform 1 0 41552 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_423
timestamp 1669390400
transform 1 0 48720 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_487
timestamp 1669390400
transform 1 0 55888 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_551
timestamp 1669390400
transform 1 0 63056 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_615
timestamp 1669390400
transform 1 0 70224 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_679
timestamp 1669390400
transform 1 0 77392 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_687
timestamp 1669390400
transform 1 0 78288 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_2
timestamp 1669390400
transform 1 0 1568 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_66
timestamp 1669390400
transform 1 0 8736 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_130
timestamp 1669390400
transform 1 0 15904 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_162
timestamp 1669390400
transform 1 0 19488 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_180
timestamp 1669390400
transform 1 0 21504 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_244
timestamp 1669390400
transform 1 0 28672 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_308
timestamp 1669390400
transform 1 0 35840 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_372
timestamp 1669390400
transform 1 0 43008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_436
timestamp 1669390400
transform 1 0 50176 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_500
timestamp 1669390400
transform 1 0 57344 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_532
timestamp 1669390400
transform 1 0 60928 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_534
timestamp 1669390400
transform 1 0 61152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_537
timestamp 1669390400
transform 1 0 61488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_601
timestamp 1669390400
transform 1 0 68656 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_665
timestamp 1669390400
transform 1 0 75824 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_681
timestamp 1669390400
transform 1 0 77616 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_685
timestamp 1669390400
transform 1 0 78064 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_687
timestamp 1669390400
transform 1 0 78288 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1669390400
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_66
timestamp 1669390400
transform 1 0 8736 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_130
timestamp 1669390400
transform 1 0 15904 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_194
timestamp 1669390400
transform 1 0 23072 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_258
timestamp 1669390400
transform 1 0 30240 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_322
timestamp 1669390400
transform 1 0 37408 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_354
timestamp 1669390400
transform 1 0 40992 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_356
timestamp 1669390400
transform 1 0 41216 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_359
timestamp 1669390400
transform 1 0 41552 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_423
timestamp 1669390400
transform 1 0 48720 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_487
timestamp 1669390400
transform 1 0 55888 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_551
timestamp 1669390400
transform 1 0 63056 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_615
timestamp 1669390400
transform 1 0 70224 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_679
timestamp 1669390400
transform 1 0 77392 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_687
timestamp 1669390400
transform 1 0 78288 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_2
timestamp 1669390400
transform 1 0 1568 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_66
timestamp 1669390400
transform 1 0 8736 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_130
timestamp 1669390400
transform 1 0 15904 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_162
timestamp 1669390400
transform 1 0 19488 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_180
timestamp 1669390400
transform 1 0 21504 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_244
timestamp 1669390400
transform 1 0 28672 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_308
timestamp 1669390400
transform 1 0 35840 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_372
timestamp 1669390400
transform 1 0 43008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_436
timestamp 1669390400
transform 1 0 50176 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_500
timestamp 1669390400
transform 1 0 57344 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_532
timestamp 1669390400
transform 1 0 60928 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_534
timestamp 1669390400
transform 1 0 61152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_537
timestamp 1669390400
transform 1 0 61488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_601
timestamp 1669390400
transform 1 0 68656 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_665
timestamp 1669390400
transform 1 0 75824 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_681
timestamp 1669390400
transform 1 0 77616 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_685
timestamp 1669390400
transform 1 0 78064 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_687
timestamp 1669390400
transform 1 0 78288 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_2
timestamp 1669390400
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_66
timestamp 1669390400
transform 1 0 8736 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_130
timestamp 1669390400
transform 1 0 15904 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_194
timestamp 1669390400
transform 1 0 23072 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_258
timestamp 1669390400
transform 1 0 30240 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_322
timestamp 1669390400
transform 1 0 37408 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_354
timestamp 1669390400
transform 1 0 40992 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_356
timestamp 1669390400
transform 1 0 41216 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_359
timestamp 1669390400
transform 1 0 41552 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_423
timestamp 1669390400
transform 1 0 48720 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_487
timestamp 1669390400
transform 1 0 55888 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_551
timestamp 1669390400
transform 1 0 63056 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_615
timestamp 1669390400
transform 1 0 70224 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_679
timestamp 1669390400
transform 1 0 77392 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_687
timestamp 1669390400
transform 1 0 78288 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_2
timestamp 1669390400
transform 1 0 1568 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_66
timestamp 1669390400
transform 1 0 8736 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_130
timestamp 1669390400
transform 1 0 15904 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_162
timestamp 1669390400
transform 1 0 19488 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_180
timestamp 1669390400
transform 1 0 21504 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_244
timestamp 1669390400
transform 1 0 28672 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_308
timestamp 1669390400
transform 1 0 35840 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_372
timestamp 1669390400
transform 1 0 43008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_436
timestamp 1669390400
transform 1 0 50176 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_500
timestamp 1669390400
transform 1 0 57344 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_532
timestamp 1669390400
transform 1 0 60928 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_534
timestamp 1669390400
transform 1 0 61152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_537
timestamp 1669390400
transform 1 0 61488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_601
timestamp 1669390400
transform 1 0 68656 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_665
timestamp 1669390400
transform 1 0 75824 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_681
timestamp 1669390400
transform 1 0 77616 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_685
timestamp 1669390400
transform 1 0 78064 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_687
timestamp 1669390400
transform 1 0 78288 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1669390400
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_66
timestamp 1669390400
transform 1 0 8736 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_130
timestamp 1669390400
transform 1 0 15904 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_194
timestamp 1669390400
transform 1 0 23072 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_258
timestamp 1669390400
transform 1 0 30240 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_322
timestamp 1669390400
transform 1 0 37408 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_354
timestamp 1669390400
transform 1 0 40992 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_356
timestamp 1669390400
transform 1 0 41216 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_359
timestamp 1669390400
transform 1 0 41552 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_423
timestamp 1669390400
transform 1 0 48720 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_487
timestamp 1669390400
transform 1 0 55888 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_551
timestamp 1669390400
transform 1 0 63056 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_615
timestamp 1669390400
transform 1 0 70224 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_679
timestamp 1669390400
transform 1 0 77392 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_687
timestamp 1669390400
transform 1 0 78288 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_2
timestamp 1669390400
transform 1 0 1568 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_66
timestamp 1669390400
transform 1 0 8736 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_130
timestamp 1669390400
transform 1 0 15904 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_162
timestamp 1669390400
transform 1 0 19488 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_180
timestamp 1669390400
transform 1 0 21504 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_244
timestamp 1669390400
transform 1 0 28672 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_308
timestamp 1669390400
transform 1 0 35840 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_372
timestamp 1669390400
transform 1 0 43008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_436
timestamp 1669390400
transform 1 0 50176 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_500
timestamp 1669390400
transform 1 0 57344 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_532
timestamp 1669390400
transform 1 0 60928 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_534
timestamp 1669390400
transform 1 0 61152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_537
timestamp 1669390400
transform 1 0 61488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_601
timestamp 1669390400
transform 1 0 68656 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_665
timestamp 1669390400
transform 1 0 75824 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_681
timestamp 1669390400
transform 1 0 77616 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_685
timestamp 1669390400
transform 1 0 78064 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_687
timestamp 1669390400
transform 1 0 78288 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1669390400
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_66
timestamp 1669390400
transform 1 0 8736 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_130
timestamp 1669390400
transform 1 0 15904 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_194
timestamp 1669390400
transform 1 0 23072 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_258
timestamp 1669390400
transform 1 0 30240 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_322
timestamp 1669390400
transform 1 0 37408 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_354
timestamp 1669390400
transform 1 0 40992 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_356
timestamp 1669390400
transform 1 0 41216 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_359
timestamp 1669390400
transform 1 0 41552 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_423
timestamp 1669390400
transform 1 0 48720 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_487
timestamp 1669390400
transform 1 0 55888 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_551
timestamp 1669390400
transform 1 0 63056 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_615
timestamp 1669390400
transform 1 0 70224 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_679
timestamp 1669390400
transform 1 0 77392 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_687
timestamp 1669390400
transform 1 0 78288 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_2
timestamp 1669390400
transform 1 0 1568 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_66
timestamp 1669390400
transform 1 0 8736 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_130
timestamp 1669390400
transform 1 0 15904 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_162
timestamp 1669390400
transform 1 0 19488 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_180
timestamp 1669390400
transform 1 0 21504 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_244
timestamp 1669390400
transform 1 0 28672 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_308
timestamp 1669390400
transform 1 0 35840 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_372
timestamp 1669390400
transform 1 0 43008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_436
timestamp 1669390400
transform 1 0 50176 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_500
timestamp 1669390400
transform 1 0 57344 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_532
timestamp 1669390400
transform 1 0 60928 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_534
timestamp 1669390400
transform 1 0 61152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_537
timestamp 1669390400
transform 1 0 61488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_601
timestamp 1669390400
transform 1 0 68656 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_665
timestamp 1669390400
transform 1 0 75824 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_681
timestamp 1669390400
transform 1 0 77616 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_685
timestamp 1669390400
transform 1 0 78064 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_687
timestamp 1669390400
transform 1 0 78288 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1669390400
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_66
timestamp 1669390400
transform 1 0 8736 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_130
timestamp 1669390400
transform 1 0 15904 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_194
timestamp 1669390400
transform 1 0 23072 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_258
timestamp 1669390400
transform 1 0 30240 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_322
timestamp 1669390400
transform 1 0 37408 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_354
timestamp 1669390400
transform 1 0 40992 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_356
timestamp 1669390400
transform 1 0 41216 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_359
timestamp 1669390400
transform 1 0 41552 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_423
timestamp 1669390400
transform 1 0 48720 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_487
timestamp 1669390400
transform 1 0 55888 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_551
timestamp 1669390400
transform 1 0 63056 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_615
timestamp 1669390400
transform 1 0 70224 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_679
timestamp 1669390400
transform 1 0 77392 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_687
timestamp 1669390400
transform 1 0 78288 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_2
timestamp 1669390400
transform 1 0 1568 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_66
timestamp 1669390400
transform 1 0 8736 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_130
timestamp 1669390400
transform 1 0 15904 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_162
timestamp 1669390400
transform 1 0 19488 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_180
timestamp 1669390400
transform 1 0 21504 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_244
timestamp 1669390400
transform 1 0 28672 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_308
timestamp 1669390400
transform 1 0 35840 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_372
timestamp 1669390400
transform 1 0 43008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_436
timestamp 1669390400
transform 1 0 50176 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_500
timestamp 1669390400
transform 1 0 57344 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_532
timestamp 1669390400
transform 1 0 60928 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_534
timestamp 1669390400
transform 1 0 61152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_537
timestamp 1669390400
transform 1 0 61488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_601
timestamp 1669390400
transform 1 0 68656 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_665
timestamp 1669390400
transform 1 0 75824 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_681
timestamp 1669390400
transform 1 0 77616 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_685
timestamp 1669390400
transform 1 0 78064 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_687
timestamp 1669390400
transform 1 0 78288 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1669390400
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_66
timestamp 1669390400
transform 1 0 8736 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_130
timestamp 1669390400
transform 1 0 15904 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_194
timestamp 1669390400
transform 1 0 23072 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_258
timestamp 1669390400
transform 1 0 30240 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_322
timestamp 1669390400
transform 1 0 37408 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_354
timestamp 1669390400
transform 1 0 40992 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_356
timestamp 1669390400
transform 1 0 41216 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_359
timestamp 1669390400
transform 1 0 41552 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_423
timestamp 1669390400
transform 1 0 48720 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_487
timestamp 1669390400
transform 1 0 55888 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_551
timestamp 1669390400
transform 1 0 63056 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_615
timestamp 1669390400
transform 1 0 70224 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_679
timestamp 1669390400
transform 1 0 77392 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_687
timestamp 1669390400
transform 1 0 78288 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_2
timestamp 1669390400
transform 1 0 1568 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_66
timestamp 1669390400
transform 1 0 8736 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_130
timestamp 1669390400
transform 1 0 15904 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_162
timestamp 1669390400
transform 1 0 19488 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_180
timestamp 1669390400
transform 1 0 21504 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_244
timestamp 1669390400
transform 1 0 28672 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_308
timestamp 1669390400
transform 1 0 35840 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_372
timestamp 1669390400
transform 1 0 43008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_436
timestamp 1669390400
transform 1 0 50176 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_500
timestamp 1669390400
transform 1 0 57344 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_532
timestamp 1669390400
transform 1 0 60928 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_534
timestamp 1669390400
transform 1 0 61152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_537
timestamp 1669390400
transform 1 0 61488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_601
timestamp 1669390400
transform 1 0 68656 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_665
timestamp 1669390400
transform 1 0 75824 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_681
timestamp 1669390400
transform 1 0 77616 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_685
timestamp 1669390400
transform 1 0 78064 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_687
timestamp 1669390400
transform 1 0 78288 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_2
timestamp 1669390400
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_66
timestamp 1669390400
transform 1 0 8736 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_130
timestamp 1669390400
transform 1 0 15904 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_194
timestamp 1669390400
transform 1 0 23072 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_258
timestamp 1669390400
transform 1 0 30240 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_322
timestamp 1669390400
transform 1 0 37408 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_354
timestamp 1669390400
transform 1 0 40992 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_356
timestamp 1669390400
transform 1 0 41216 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_359
timestamp 1669390400
transform 1 0 41552 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_423
timestamp 1669390400
transform 1 0 48720 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_487
timestamp 1669390400
transform 1 0 55888 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_551
timestamp 1669390400
transform 1 0 63056 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_615
timestamp 1669390400
transform 1 0 70224 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_679
timestamp 1669390400
transform 1 0 77392 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_687
timestamp 1669390400
transform 1 0 78288 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_2
timestamp 1669390400
transform 1 0 1568 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_66
timestamp 1669390400
transform 1 0 8736 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_130
timestamp 1669390400
transform 1 0 15904 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_162
timestamp 1669390400
transform 1 0 19488 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_180
timestamp 1669390400
transform 1 0 21504 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_244
timestamp 1669390400
transform 1 0 28672 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_308
timestamp 1669390400
transform 1 0 35840 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_372
timestamp 1669390400
transform 1 0 43008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_436
timestamp 1669390400
transform 1 0 50176 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_500
timestamp 1669390400
transform 1 0 57344 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_532
timestamp 1669390400
transform 1 0 60928 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_534
timestamp 1669390400
transform 1 0 61152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_537
timestamp 1669390400
transform 1 0 61488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_601
timestamp 1669390400
transform 1 0 68656 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_665
timestamp 1669390400
transform 1 0 75824 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_681
timestamp 1669390400
transform 1 0 77616 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_685
timestamp 1669390400
transform 1 0 78064 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_687
timestamp 1669390400
transform 1 0 78288 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_2
timestamp 1669390400
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_66
timestamp 1669390400
transform 1 0 8736 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_130
timestamp 1669390400
transform 1 0 15904 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_194
timestamp 1669390400
transform 1 0 23072 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_258
timestamp 1669390400
transform 1 0 30240 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_322
timestamp 1669390400
transform 1 0 37408 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_354
timestamp 1669390400
transform 1 0 40992 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_356
timestamp 1669390400
transform 1 0 41216 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_359
timestamp 1669390400
transform 1 0 41552 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_423
timestamp 1669390400
transform 1 0 48720 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_487
timestamp 1669390400
transform 1 0 55888 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_551
timestamp 1669390400
transform 1 0 63056 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_615
timestamp 1669390400
transform 1 0 70224 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_679
timestamp 1669390400
transform 1 0 77392 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_687
timestamp 1669390400
transform 1 0 78288 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_2
timestamp 1669390400
transform 1 0 1568 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_66
timestamp 1669390400
transform 1 0 8736 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_130
timestamp 1669390400
transform 1 0 15904 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_162
timestamp 1669390400
transform 1 0 19488 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_180
timestamp 1669390400
transform 1 0 21504 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_244
timestamp 1669390400
transform 1 0 28672 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_308
timestamp 1669390400
transform 1 0 35840 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_372
timestamp 1669390400
transform 1 0 43008 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_436
timestamp 1669390400
transform 1 0 50176 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_500
timestamp 1669390400
transform 1 0 57344 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_532
timestamp 1669390400
transform 1 0 60928 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_534
timestamp 1669390400
transform 1 0 61152 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_537
timestamp 1669390400
transform 1 0 61488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_601
timestamp 1669390400
transform 1 0 68656 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_665
timestamp 1669390400
transform 1 0 75824 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_681
timestamp 1669390400
transform 1 0 77616 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_685
timestamp 1669390400
transform 1 0 78064 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_687
timestamp 1669390400
transform 1 0 78288 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_2
timestamp 1669390400
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_66
timestamp 1669390400
transform 1 0 8736 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_130
timestamp 1669390400
transform 1 0 15904 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_194
timestamp 1669390400
transform 1 0 23072 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_258
timestamp 1669390400
transform 1 0 30240 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_322
timestamp 1669390400
transform 1 0 37408 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_354
timestamp 1669390400
transform 1 0 40992 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_356
timestamp 1669390400
transform 1 0 41216 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_359
timestamp 1669390400
transform 1 0 41552 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_423
timestamp 1669390400
transform 1 0 48720 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_487
timestamp 1669390400
transform 1 0 55888 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_551
timestamp 1669390400
transform 1 0 63056 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_615
timestamp 1669390400
transform 1 0 70224 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_679
timestamp 1669390400
transform 1 0 77392 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_687
timestamp 1669390400
transform 1 0 78288 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_2
timestamp 1669390400
transform 1 0 1568 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_66
timestamp 1669390400
transform 1 0 8736 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_130
timestamp 1669390400
transform 1 0 15904 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_162
timestamp 1669390400
transform 1 0 19488 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_180
timestamp 1669390400
transform 1 0 21504 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_244
timestamp 1669390400
transform 1 0 28672 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_308
timestamp 1669390400
transform 1 0 35840 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_372
timestamp 1669390400
transform 1 0 43008 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_436
timestamp 1669390400
transform 1 0 50176 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_500
timestamp 1669390400
transform 1 0 57344 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_532
timestamp 1669390400
transform 1 0 60928 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_534
timestamp 1669390400
transform 1 0 61152 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_537
timestamp 1669390400
transform 1 0 61488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_46_601
timestamp 1669390400
transform 1 0 68656 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_665
timestamp 1669390400
transform 1 0 75824 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_681
timestamp 1669390400
transform 1 0 77616 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_685
timestamp 1669390400
transform 1 0 78064 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_687
timestamp 1669390400
transform 1 0 78288 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_2
timestamp 1669390400
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_66
timestamp 1669390400
transform 1 0 8736 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_130
timestamp 1669390400
transform 1 0 15904 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_194
timestamp 1669390400
transform 1 0 23072 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_258
timestamp 1669390400
transform 1 0 30240 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_322
timestamp 1669390400
transform 1 0 37408 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_354
timestamp 1669390400
transform 1 0 40992 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_356
timestamp 1669390400
transform 1 0 41216 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_359
timestamp 1669390400
transform 1 0 41552 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_423
timestamp 1669390400
transform 1 0 48720 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_487
timestamp 1669390400
transform 1 0 55888 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_551
timestamp 1669390400
transform 1 0 63056 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_615
timestamp 1669390400
transform 1 0 70224 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_679
timestamp 1669390400
transform 1 0 77392 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_687
timestamp 1669390400
transform 1 0 78288 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_2
timestamp 1669390400
transform 1 0 1568 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_66
timestamp 1669390400
transform 1 0 8736 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_130
timestamp 1669390400
transform 1 0 15904 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_162
timestamp 1669390400
transform 1 0 19488 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_180
timestamp 1669390400
transform 1 0 21504 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_244
timestamp 1669390400
transform 1 0 28672 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_308
timestamp 1669390400
transform 1 0 35840 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_372
timestamp 1669390400
transform 1 0 43008 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_436
timestamp 1669390400
transform 1 0 50176 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_500
timestamp 1669390400
transform 1 0 57344 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_532
timestamp 1669390400
transform 1 0 60928 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_534
timestamp 1669390400
transform 1 0 61152 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_537
timestamp 1669390400
transform 1 0 61488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_48_601
timestamp 1669390400
transform 1 0 68656 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_665
timestamp 1669390400
transform 1 0 75824 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_681
timestamp 1669390400
transform 1 0 77616 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_685
timestamp 1669390400
transform 1 0 78064 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_687
timestamp 1669390400
transform 1 0 78288 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_2
timestamp 1669390400
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_66
timestamp 1669390400
transform 1 0 8736 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_130
timestamp 1669390400
transform 1 0 15904 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_194
timestamp 1669390400
transform 1 0 23072 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_258
timestamp 1669390400
transform 1 0 30240 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_322
timestamp 1669390400
transform 1 0 37408 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_354
timestamp 1669390400
transform 1 0 40992 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_356
timestamp 1669390400
transform 1 0 41216 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_359
timestamp 1669390400
transform 1 0 41552 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_423
timestamp 1669390400
transform 1 0 48720 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_487
timestamp 1669390400
transform 1 0 55888 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_551
timestamp 1669390400
transform 1 0 63056 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_615
timestamp 1669390400
transform 1 0 70224 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_679
timestamp 1669390400
transform 1 0 77392 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_687
timestamp 1669390400
transform 1 0 78288 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_2
timestamp 1669390400
transform 1 0 1568 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_66
timestamp 1669390400
transform 1 0 8736 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_130
timestamp 1669390400
transform 1 0 15904 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_162
timestamp 1669390400
transform 1 0 19488 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_180
timestamp 1669390400
transform 1 0 21504 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_244
timestamp 1669390400
transform 1 0 28672 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_308
timestamp 1669390400
transform 1 0 35840 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_372
timestamp 1669390400
transform 1 0 43008 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_436
timestamp 1669390400
transform 1 0 50176 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_500
timestamp 1669390400
transform 1 0 57344 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_532
timestamp 1669390400
transform 1 0 60928 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_534
timestamp 1669390400
transform 1 0 61152 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_537
timestamp 1669390400
transform 1 0 61488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_601
timestamp 1669390400
transform 1 0 68656 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_665
timestamp 1669390400
transform 1 0 75824 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_681
timestamp 1669390400
transform 1 0 77616 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_685
timestamp 1669390400
transform 1 0 78064 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_687
timestamp 1669390400
transform 1 0 78288 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_2
timestamp 1669390400
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_66
timestamp 1669390400
transform 1 0 8736 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_130
timestamp 1669390400
transform 1 0 15904 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_194
timestamp 1669390400
transform 1 0 23072 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_258
timestamp 1669390400
transform 1 0 30240 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_322
timestamp 1669390400
transform 1 0 37408 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_354
timestamp 1669390400
transform 1 0 40992 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_356
timestamp 1669390400
transform 1 0 41216 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_359
timestamp 1669390400
transform 1 0 41552 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_423
timestamp 1669390400
transform 1 0 48720 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_487
timestamp 1669390400
transform 1 0 55888 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_551
timestamp 1669390400
transform 1 0 63056 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_615
timestamp 1669390400
transform 1 0 70224 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_679
timestamp 1669390400
transform 1 0 77392 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_687
timestamp 1669390400
transform 1 0 78288 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_2
timestamp 1669390400
transform 1 0 1568 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_66
timestamp 1669390400
transform 1 0 8736 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_130
timestamp 1669390400
transform 1 0 15904 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_162
timestamp 1669390400
transform 1 0 19488 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_180
timestamp 1669390400
transform 1 0 21504 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_244
timestamp 1669390400
transform 1 0 28672 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_308
timestamp 1669390400
transform 1 0 35840 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_372
timestamp 1669390400
transform 1 0 43008 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_436
timestamp 1669390400
transform 1 0 50176 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_500
timestamp 1669390400
transform 1 0 57344 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_532
timestamp 1669390400
transform 1 0 60928 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_534
timestamp 1669390400
transform 1 0 61152 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_537
timestamp 1669390400
transform 1 0 61488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_52_601
timestamp 1669390400
transform 1 0 68656 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_665
timestamp 1669390400
transform 1 0 75824 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_681
timestamp 1669390400
transform 1 0 77616 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_685
timestamp 1669390400
transform 1 0 78064 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_687
timestamp 1669390400
transform 1 0 78288 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_2
timestamp 1669390400
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_66
timestamp 1669390400
transform 1 0 8736 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_130
timestamp 1669390400
transform 1 0 15904 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_194
timestamp 1669390400
transform 1 0 23072 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_258
timestamp 1669390400
transform 1 0 30240 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_322
timestamp 1669390400
transform 1 0 37408 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_354
timestamp 1669390400
transform 1 0 40992 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_356
timestamp 1669390400
transform 1 0 41216 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_359
timestamp 1669390400
transform 1 0 41552 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_423
timestamp 1669390400
transform 1 0 48720 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_487
timestamp 1669390400
transform 1 0 55888 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_551
timestamp 1669390400
transform 1 0 63056 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_615
timestamp 1669390400
transform 1 0 70224 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_679
timestamp 1669390400
transform 1 0 77392 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_687
timestamp 1669390400
transform 1 0 78288 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_2
timestamp 1669390400
transform 1 0 1568 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_66
timestamp 1669390400
transform 1 0 8736 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_130
timestamp 1669390400
transform 1 0 15904 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_162
timestamp 1669390400
transform 1 0 19488 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_180
timestamp 1669390400
transform 1 0 21504 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_244
timestamp 1669390400
transform 1 0 28672 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_308
timestamp 1669390400
transform 1 0 35840 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_372
timestamp 1669390400
transform 1 0 43008 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_436
timestamp 1669390400
transform 1 0 50176 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_500
timestamp 1669390400
transform 1 0 57344 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_532
timestamp 1669390400
transform 1 0 60928 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_534
timestamp 1669390400
transform 1 0 61152 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_537
timestamp 1669390400
transform 1 0 61488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_601
timestamp 1669390400
transform 1 0 68656 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_665
timestamp 1669390400
transform 1 0 75824 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_681
timestamp 1669390400
transform 1 0 77616 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_685
timestamp 1669390400
transform 1 0 78064 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_687
timestamp 1669390400
transform 1 0 78288 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_2
timestamp 1669390400
transform 1 0 1568 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_66
timestamp 1669390400
transform 1 0 8736 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_130
timestamp 1669390400
transform 1 0 15904 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_194
timestamp 1669390400
transform 1 0 23072 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_258
timestamp 1669390400
transform 1 0 30240 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_322
timestamp 1669390400
transform 1 0 37408 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_354
timestamp 1669390400
transform 1 0 40992 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_356
timestamp 1669390400
transform 1 0 41216 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_359
timestamp 1669390400
transform 1 0 41552 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_423
timestamp 1669390400
transform 1 0 48720 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_487
timestamp 1669390400
transform 1 0 55888 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_551
timestamp 1669390400
transform 1 0 63056 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_615
timestamp 1669390400
transform 1 0 70224 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_679
timestamp 1669390400
transform 1 0 77392 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_687
timestamp 1669390400
transform 1 0 78288 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_2
timestamp 1669390400
transform 1 0 1568 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_66
timestamp 1669390400
transform 1 0 8736 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_130
timestamp 1669390400
transform 1 0 15904 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_162
timestamp 1669390400
transform 1 0 19488 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_180
timestamp 1669390400
transform 1 0 21504 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_244
timestamp 1669390400
transform 1 0 28672 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_308
timestamp 1669390400
transform 1 0 35840 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_372
timestamp 1669390400
transform 1 0 43008 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_436
timestamp 1669390400
transform 1 0 50176 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_500
timestamp 1669390400
transform 1 0 57344 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_532
timestamp 1669390400
transform 1 0 60928 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_534
timestamp 1669390400
transform 1 0 61152 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_537
timestamp 1669390400
transform 1 0 61488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_56_601
timestamp 1669390400
transform 1 0 68656 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_665
timestamp 1669390400
transform 1 0 75824 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_681
timestamp 1669390400
transform 1 0 77616 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_685
timestamp 1669390400
transform 1 0 78064 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_687
timestamp 1669390400
transform 1 0 78288 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_2
timestamp 1669390400
transform 1 0 1568 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_66
timestamp 1669390400
transform 1 0 8736 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_130
timestamp 1669390400
transform 1 0 15904 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_194
timestamp 1669390400
transform 1 0 23072 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_258
timestamp 1669390400
transform 1 0 30240 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_322
timestamp 1669390400
transform 1 0 37408 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_354
timestamp 1669390400
transform 1 0 40992 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_356
timestamp 1669390400
transform 1 0 41216 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_359
timestamp 1669390400
transform 1 0 41552 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_423
timestamp 1669390400
transform 1 0 48720 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_487
timestamp 1669390400
transform 1 0 55888 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_551
timestamp 1669390400
transform 1 0 63056 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_615
timestamp 1669390400
transform 1 0 70224 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_679
timestamp 1669390400
transform 1 0 77392 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_687
timestamp 1669390400
transform 1 0 78288 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_2
timestamp 1669390400
transform 1 0 1568 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_66
timestamp 1669390400
transform 1 0 8736 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_130
timestamp 1669390400
transform 1 0 15904 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_162
timestamp 1669390400
transform 1 0 19488 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_180
timestamp 1669390400
transform 1 0 21504 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_244
timestamp 1669390400
transform 1 0 28672 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_308
timestamp 1669390400
transform 1 0 35840 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_372
timestamp 1669390400
transform 1 0 43008 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_436
timestamp 1669390400
transform 1 0 50176 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_500
timestamp 1669390400
transform 1 0 57344 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_532
timestamp 1669390400
transform 1 0 60928 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_534
timestamp 1669390400
transform 1 0 61152 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_537
timestamp 1669390400
transform 1 0 61488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_58_601
timestamp 1669390400
transform 1 0 68656 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_665
timestamp 1669390400
transform 1 0 75824 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_681
timestamp 1669390400
transform 1 0 77616 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_685
timestamp 1669390400
transform 1 0 78064 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_687
timestamp 1669390400
transform 1 0 78288 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_2
timestamp 1669390400
transform 1 0 1568 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_66
timestamp 1669390400
transform 1 0 8736 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_130
timestamp 1669390400
transform 1 0 15904 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_194
timestamp 1669390400
transform 1 0 23072 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_258
timestamp 1669390400
transform 1 0 30240 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_59_322
timestamp 1669390400
transform 1 0 37408 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_354
timestamp 1669390400
transform 1 0 40992 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_356
timestamp 1669390400
transform 1 0 41216 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_359
timestamp 1669390400
transform 1 0 41552 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_423
timestamp 1669390400
transform 1 0 48720 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_487
timestamp 1669390400
transform 1 0 55888 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_551
timestamp 1669390400
transform 1 0 63056 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_615
timestamp 1669390400
transform 1 0 70224 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_679
timestamp 1669390400
transform 1 0 77392 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_687
timestamp 1669390400
transform 1 0 78288 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_2
timestamp 1669390400
transform 1 0 1568 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_66
timestamp 1669390400
transform 1 0 8736 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_130
timestamp 1669390400
transform 1 0 15904 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_162
timestamp 1669390400
transform 1 0 19488 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_180
timestamp 1669390400
transform 1 0 21504 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_244
timestamp 1669390400
transform 1 0 28672 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_308
timestamp 1669390400
transform 1 0 35840 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_372
timestamp 1669390400
transform 1 0 43008 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_436
timestamp 1669390400
transform 1 0 50176 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_500
timestamp 1669390400
transform 1 0 57344 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_532
timestamp 1669390400
transform 1 0 60928 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_534
timestamp 1669390400
transform 1 0 61152 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_537
timestamp 1669390400
transform 1 0 61488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_601
timestamp 1669390400
transform 1 0 68656 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_665
timestamp 1669390400
transform 1 0 75824 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_681
timestamp 1669390400
transform 1 0 77616 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_685
timestamp 1669390400
transform 1 0 78064 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_687
timestamp 1669390400
transform 1 0 78288 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_2
timestamp 1669390400
transform 1 0 1568 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_66
timestamp 1669390400
transform 1 0 8736 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_130
timestamp 1669390400
transform 1 0 15904 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_194
timestamp 1669390400
transform 1 0 23072 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_258
timestamp 1669390400
transform 1 0 30240 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_322
timestamp 1669390400
transform 1 0 37408 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_354
timestamp 1669390400
transform 1 0 40992 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_356
timestamp 1669390400
transform 1 0 41216 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_359
timestamp 1669390400
transform 1 0 41552 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_423
timestamp 1669390400
transform 1 0 48720 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_487
timestamp 1669390400
transform 1 0 55888 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_551
timestamp 1669390400
transform 1 0 63056 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_615
timestamp 1669390400
transform 1 0 70224 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_679
timestamp 1669390400
transform 1 0 77392 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_687
timestamp 1669390400
transform 1 0 78288 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_2
timestamp 1669390400
transform 1 0 1568 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_66
timestamp 1669390400
transform 1 0 8736 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_130
timestamp 1669390400
transform 1 0 15904 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_162
timestamp 1669390400
transform 1 0 19488 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_180
timestamp 1669390400
transform 1 0 21504 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_244
timestamp 1669390400
transform 1 0 28672 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_308
timestamp 1669390400
transform 1 0 35840 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_372
timestamp 1669390400
transform 1 0 43008 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_436
timestamp 1669390400
transform 1 0 50176 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_500
timestamp 1669390400
transform 1 0 57344 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_532
timestamp 1669390400
transform 1 0 60928 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_534
timestamp 1669390400
transform 1 0 61152 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_537
timestamp 1669390400
transform 1 0 61488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_601
timestamp 1669390400
transform 1 0 68656 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_665
timestamp 1669390400
transform 1 0 75824 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_681
timestamp 1669390400
transform 1 0 77616 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_685
timestamp 1669390400
transform 1 0 78064 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_687
timestamp 1669390400
transform 1 0 78288 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_2
timestamp 1669390400
transform 1 0 1568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_66
timestamp 1669390400
transform 1 0 8736 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_130
timestamp 1669390400
transform 1 0 15904 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_194
timestamp 1669390400
transform 1 0 23072 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_258
timestamp 1669390400
transform 1 0 30240 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_63_322
timestamp 1669390400
transform 1 0 37408 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_354
timestamp 1669390400
transform 1 0 40992 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_356
timestamp 1669390400
transform 1 0 41216 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_359
timestamp 1669390400
transform 1 0 41552 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_423
timestamp 1669390400
transform 1 0 48720 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_487
timestamp 1669390400
transform 1 0 55888 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_551
timestamp 1669390400
transform 1 0 63056 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_615
timestamp 1669390400
transform 1 0 70224 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_679
timestamp 1669390400
transform 1 0 77392 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_687
timestamp 1669390400
transform 1 0 78288 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_2
timestamp 1669390400
transform 1 0 1568 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_66
timestamp 1669390400
transform 1 0 8736 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_130
timestamp 1669390400
transform 1 0 15904 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_162
timestamp 1669390400
transform 1 0 19488 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_180
timestamp 1669390400
transform 1 0 21504 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_244
timestamp 1669390400
transform 1 0 28672 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_308
timestamp 1669390400
transform 1 0 35840 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_372
timestamp 1669390400
transform 1 0 43008 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_436
timestamp 1669390400
transform 1 0 50176 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_500
timestamp 1669390400
transform 1 0 57344 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_532
timestamp 1669390400
transform 1 0 60928 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_534
timestamp 1669390400
transform 1 0 61152 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_537
timestamp 1669390400
transform 1 0 61488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_601
timestamp 1669390400
transform 1 0 68656 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_665
timestamp 1669390400
transform 1 0 75824 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_681
timestamp 1669390400
transform 1 0 77616 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_685
timestamp 1669390400
transform 1 0 78064 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_687
timestamp 1669390400
transform 1 0 78288 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_2
timestamp 1669390400
transform 1 0 1568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_66
timestamp 1669390400
transform 1 0 8736 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_130
timestamp 1669390400
transform 1 0 15904 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_194
timestamp 1669390400
transform 1 0 23072 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_258
timestamp 1669390400
transform 1 0 30240 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_322
timestamp 1669390400
transform 1 0 37408 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_354
timestamp 1669390400
transform 1 0 40992 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_356
timestamp 1669390400
transform 1 0 41216 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_359
timestamp 1669390400
transform 1 0 41552 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_423
timestamp 1669390400
transform 1 0 48720 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_487
timestamp 1669390400
transform 1 0 55888 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_551
timestamp 1669390400
transform 1 0 63056 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_615
timestamp 1669390400
transform 1 0 70224 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_679
timestamp 1669390400
transform 1 0 77392 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_687
timestamp 1669390400
transform 1 0 78288 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_2
timestamp 1669390400
transform 1 0 1568 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_66
timestamp 1669390400
transform 1 0 8736 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_130
timestamp 1669390400
transform 1 0 15904 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_162
timestamp 1669390400
transform 1 0 19488 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_180
timestamp 1669390400
transform 1 0 21504 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_244
timestamp 1669390400
transform 1 0 28672 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_308
timestamp 1669390400
transform 1 0 35840 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_372
timestamp 1669390400
transform 1 0 43008 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_436
timestamp 1669390400
transform 1 0 50176 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_500
timestamp 1669390400
transform 1 0 57344 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_532
timestamp 1669390400
transform 1 0 60928 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_534
timestamp 1669390400
transform 1 0 61152 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_537
timestamp 1669390400
transform 1 0 61488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_601
timestamp 1669390400
transform 1 0 68656 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_665
timestamp 1669390400
transform 1 0 75824 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_681
timestamp 1669390400
transform 1 0 77616 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_685
timestamp 1669390400
transform 1 0 78064 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_687
timestamp 1669390400
transform 1 0 78288 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_2
timestamp 1669390400
transform 1 0 1568 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_66
timestamp 1669390400
transform 1 0 8736 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_130
timestamp 1669390400
transform 1 0 15904 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_194
timestamp 1669390400
transform 1 0 23072 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_258
timestamp 1669390400
transform 1 0 30240 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_322
timestamp 1669390400
transform 1 0 37408 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_354
timestamp 1669390400
transform 1 0 40992 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_356
timestamp 1669390400
transform 1 0 41216 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_359
timestamp 1669390400
transform 1 0 41552 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_423
timestamp 1669390400
transform 1 0 48720 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_487
timestamp 1669390400
transform 1 0 55888 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_551
timestamp 1669390400
transform 1 0 63056 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_67_615
timestamp 1669390400
transform 1 0 70224 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_679
timestamp 1669390400
transform 1 0 77392 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_687
timestamp 1669390400
transform 1 0 78288 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_2
timestamp 1669390400
transform 1 0 1568 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_66
timestamp 1669390400
transform 1 0 8736 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_68_130
timestamp 1669390400
transform 1 0 15904 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_162
timestamp 1669390400
transform 1 0 19488 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_180
timestamp 1669390400
transform 1 0 21504 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_244
timestamp 1669390400
transform 1 0 28672 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_308
timestamp 1669390400
transform 1 0 35840 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_372
timestamp 1669390400
transform 1 0 43008 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_436
timestamp 1669390400
transform 1 0 50176 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_68_500
timestamp 1669390400
transform 1 0 57344 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_532
timestamp 1669390400
transform 1 0 60928 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_534
timestamp 1669390400
transform 1 0 61152 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_537
timestamp 1669390400
transform 1 0 61488 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_68_601
timestamp 1669390400
transform 1 0 68656 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_68_665
timestamp 1669390400
transform 1 0 75824 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_68_681
timestamp 1669390400
transform 1 0 77616 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_68_685
timestamp 1669390400
transform 1 0 78064 0 1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_68_687
timestamp 1669390400
transform 1 0 78288 0 1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_2
timestamp 1669390400
transform 1 0 1568 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_66
timestamp 1669390400
transform 1 0 8736 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_130
timestamp 1669390400
transform 1 0 15904 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_194
timestamp 1669390400
transform 1 0 23072 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_258
timestamp 1669390400
transform 1 0 30240 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_69_322
timestamp 1669390400
transform 1 0 37408 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_69_354
timestamp 1669390400
transform 1 0 40992 0 -1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_356
timestamp 1669390400
transform 1 0 41216 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_359
timestamp 1669390400
transform 1 0 41552 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_423
timestamp 1669390400
transform 1 0 48720 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_487
timestamp 1669390400
transform 1 0 55888 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_551
timestamp 1669390400
transform 1 0 63056 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_69_615
timestamp 1669390400
transform 1 0 70224 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_69_679
timestamp 1669390400
transform 1 0 77392 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_69_687
timestamp 1669390400
transform 1 0 78288 0 -1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_2
timestamp 1669390400
transform 1 0 1568 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_66
timestamp 1669390400
transform 1 0 8736 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_70_130
timestamp 1669390400
transform 1 0 15904 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_70_162
timestamp 1669390400
transform 1 0 19488 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_180
timestamp 1669390400
transform 1 0 21504 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_244
timestamp 1669390400
transform 1 0 28672 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_308
timestamp 1669390400
transform 1 0 35840 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_372
timestamp 1669390400
transform 1 0 43008 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_436
timestamp 1669390400
transform 1 0 50176 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_70_500
timestamp 1669390400
transform 1 0 57344 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_532
timestamp 1669390400
transform 1 0 60928 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_534
timestamp 1669390400
transform 1 0 61152 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_537
timestamp 1669390400
transform 1 0 61488 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_70_601
timestamp 1669390400
transform 1 0 68656 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_70_665
timestamp 1669390400
transform 1 0 75824 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_70_681
timestamp 1669390400
transform 1 0 77616 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_70_685
timestamp 1669390400
transform 1 0 78064 0 1 58016
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_70_687
timestamp 1669390400
transform 1 0 78288 0 1 58016
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_2
timestamp 1669390400
transform 1 0 1568 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_66
timestamp 1669390400
transform 1 0 8736 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_130
timestamp 1669390400
transform 1 0 15904 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_194
timestamp 1669390400
transform 1 0 23072 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_258
timestamp 1669390400
transform 1 0 30240 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_71_322
timestamp 1669390400
transform 1 0 37408 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_71_354
timestamp 1669390400
transform 1 0 40992 0 -1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_356
timestamp 1669390400
transform 1 0 41216 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_359
timestamp 1669390400
transform 1 0 41552 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_423
timestamp 1669390400
transform 1 0 48720 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_487
timestamp 1669390400
transform 1 0 55888 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_551
timestamp 1669390400
transform 1 0 63056 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_71_615
timestamp 1669390400
transform 1 0 70224 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_71_679
timestamp 1669390400
transform 1 0 77392 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_71_687
timestamp 1669390400
transform 1 0 78288 0 -1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_2
timestamp 1669390400
transform 1 0 1568 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_66
timestamp 1669390400
transform 1 0 8736 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_72_130
timestamp 1669390400
transform 1 0 15904 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_72_162
timestamp 1669390400
transform 1 0 19488 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_180
timestamp 1669390400
transform 1 0 21504 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_244
timestamp 1669390400
transform 1 0 28672 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_308
timestamp 1669390400
transform 1 0 35840 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_372
timestamp 1669390400
transform 1 0 43008 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_436
timestamp 1669390400
transform 1 0 50176 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_72_500
timestamp 1669390400
transform 1 0 57344 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_532
timestamp 1669390400
transform 1 0 60928 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_534
timestamp 1669390400
transform 1 0 61152 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_537
timestamp 1669390400
transform 1 0 61488 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_72_601
timestamp 1669390400
transform 1 0 68656 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_72_665
timestamp 1669390400
transform 1 0 75824 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_72_681
timestamp 1669390400
transform 1 0 77616 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_72_685
timestamp 1669390400
transform 1 0 78064 0 1 59584
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_72_687
timestamp 1669390400
transform 1 0 78288 0 1 59584
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_2
timestamp 1669390400
transform 1 0 1568 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_66
timestamp 1669390400
transform 1 0 8736 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_130
timestamp 1669390400
transform 1 0 15904 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_194
timestamp 1669390400
transform 1 0 23072 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_258
timestamp 1669390400
transform 1 0 30240 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_73_322
timestamp 1669390400
transform 1 0 37408 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_73_354
timestamp 1669390400
transform 1 0 40992 0 -1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_356
timestamp 1669390400
transform 1 0 41216 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_359
timestamp 1669390400
transform 1 0 41552 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_423
timestamp 1669390400
transform 1 0 48720 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_487
timestamp 1669390400
transform 1 0 55888 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_551
timestamp 1669390400
transform 1 0 63056 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_73_615
timestamp 1669390400
transform 1 0 70224 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_73_679
timestamp 1669390400
transform 1 0 77392 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_73_687
timestamp 1669390400
transform 1 0 78288 0 -1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_2
timestamp 1669390400
transform 1 0 1568 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_66
timestamp 1669390400
transform 1 0 8736 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_74_130
timestamp 1669390400
transform 1 0 15904 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_74_162
timestamp 1669390400
transform 1 0 19488 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_180
timestamp 1669390400
transform 1 0 21504 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_244
timestamp 1669390400
transform 1 0 28672 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_308
timestamp 1669390400
transform 1 0 35840 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_372
timestamp 1669390400
transform 1 0 43008 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_436
timestamp 1669390400
transform 1 0 50176 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_74_500
timestamp 1669390400
transform 1 0 57344 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_532
timestamp 1669390400
transform 1 0 60928 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_534
timestamp 1669390400
transform 1 0 61152 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_537
timestamp 1669390400
transform 1 0 61488 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_74_601
timestamp 1669390400
transform 1 0 68656 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_74_665
timestamp 1669390400
transform 1 0 75824 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_74_681
timestamp 1669390400
transform 1 0 77616 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_74_685
timestamp 1669390400
transform 1 0 78064 0 1 61152
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_74_687
timestamp 1669390400
transform 1 0 78288 0 1 61152
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_2
timestamp 1669390400
transform 1 0 1568 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_66
timestamp 1669390400
transform 1 0 8736 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_130
timestamp 1669390400
transform 1 0 15904 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_194
timestamp 1669390400
transform 1 0 23072 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_258
timestamp 1669390400
transform 1 0 30240 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_75_322
timestamp 1669390400
transform 1 0 37408 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_75_354
timestamp 1669390400
transform 1 0 40992 0 -1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_356
timestamp 1669390400
transform 1 0 41216 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_359
timestamp 1669390400
transform 1 0 41552 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_423
timestamp 1669390400
transform 1 0 48720 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_487
timestamp 1669390400
transform 1 0 55888 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_551
timestamp 1669390400
transform 1 0 63056 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_75_615
timestamp 1669390400
transform 1 0 70224 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_75_679
timestamp 1669390400
transform 1 0 77392 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_75_687
timestamp 1669390400
transform 1 0 78288 0 -1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_2
timestamp 1669390400
transform 1 0 1568 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_66
timestamp 1669390400
transform 1 0 8736 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_76_130
timestamp 1669390400
transform 1 0 15904 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_76_162
timestamp 1669390400
transform 1 0 19488 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_180
timestamp 1669390400
transform 1 0 21504 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_244
timestamp 1669390400
transform 1 0 28672 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_308
timestamp 1669390400
transform 1 0 35840 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_372
timestamp 1669390400
transform 1 0 43008 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_436
timestamp 1669390400
transform 1 0 50176 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_76_500
timestamp 1669390400
transform 1 0 57344 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_532
timestamp 1669390400
transform 1 0 60928 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_534
timestamp 1669390400
transform 1 0 61152 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_537
timestamp 1669390400
transform 1 0 61488 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_76_601
timestamp 1669390400
transform 1 0 68656 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_76_665
timestamp 1669390400
transform 1 0 75824 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_76_681
timestamp 1669390400
transform 1 0 77616 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_76_685
timestamp 1669390400
transform 1 0 78064 0 1 62720
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_76_687
timestamp 1669390400
transform 1 0 78288 0 1 62720
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_2
timestamp 1669390400
transform 1 0 1568 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_66
timestamp 1669390400
transform 1 0 8736 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_130
timestamp 1669390400
transform 1 0 15904 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_194
timestamp 1669390400
transform 1 0 23072 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_258
timestamp 1669390400
transform 1 0 30240 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_77_322
timestamp 1669390400
transform 1 0 37408 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_77_354
timestamp 1669390400
transform 1 0 40992 0 -1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_356
timestamp 1669390400
transform 1 0 41216 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_359
timestamp 1669390400
transform 1 0 41552 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_423
timestamp 1669390400
transform 1 0 48720 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_487
timestamp 1669390400
transform 1 0 55888 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_551
timestamp 1669390400
transform 1 0 63056 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_77_615
timestamp 1669390400
transform 1 0 70224 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_77_679
timestamp 1669390400
transform 1 0 77392 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_77_687
timestamp 1669390400
transform 1 0 78288 0 -1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_2
timestamp 1669390400
transform 1 0 1568 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_66
timestamp 1669390400
transform 1 0 8736 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_78_130
timestamp 1669390400
transform 1 0 15904 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_78_162
timestamp 1669390400
transform 1 0 19488 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_180
timestamp 1669390400
transform 1 0 21504 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_244
timestamp 1669390400
transform 1 0 28672 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_308
timestamp 1669390400
transform 1 0 35840 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_372
timestamp 1669390400
transform 1 0 43008 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_436
timestamp 1669390400
transform 1 0 50176 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_78_500
timestamp 1669390400
transform 1 0 57344 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_532
timestamp 1669390400
transform 1 0 60928 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_534
timestamp 1669390400
transform 1 0 61152 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_537
timestamp 1669390400
transform 1 0 61488 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_78_601
timestamp 1669390400
transform 1 0 68656 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_78_665
timestamp 1669390400
transform 1 0 75824 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_78_681
timestamp 1669390400
transform 1 0 77616 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_78_685
timestamp 1669390400
transform 1 0 78064 0 1 64288
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_78_687
timestamp 1669390400
transform 1 0 78288 0 1 64288
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_2
timestamp 1669390400
transform 1 0 1568 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_66
timestamp 1669390400
transform 1 0 8736 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_130
timestamp 1669390400
transform 1 0 15904 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_194
timestamp 1669390400
transform 1 0 23072 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_258
timestamp 1669390400
transform 1 0 30240 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_79_322
timestamp 1669390400
transform 1 0 37408 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_79_354
timestamp 1669390400
transform 1 0 40992 0 -1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_356
timestamp 1669390400
transform 1 0 41216 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_359
timestamp 1669390400
transform 1 0 41552 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_423
timestamp 1669390400
transform 1 0 48720 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_487
timestamp 1669390400
transform 1 0 55888 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_551
timestamp 1669390400
transform 1 0 63056 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_79_615
timestamp 1669390400
transform 1 0 70224 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_79_679
timestamp 1669390400
transform 1 0 77392 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_79_687
timestamp 1669390400
transform 1 0 78288 0 -1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_2
timestamp 1669390400
transform 1 0 1568 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_66
timestamp 1669390400
transform 1 0 8736 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_130
timestamp 1669390400
transform 1 0 15904 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_80_162
timestamp 1669390400
transform 1 0 19488 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_180
timestamp 1669390400
transform 1 0 21504 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_244
timestamp 1669390400
transform 1 0 28672 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_308
timestamp 1669390400
transform 1 0 35840 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_372
timestamp 1669390400
transform 1 0 43008 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_436
timestamp 1669390400
transform 1 0 50176 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_80_500
timestamp 1669390400
transform 1 0 57344 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_532
timestamp 1669390400
transform 1 0 60928 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_534
timestamp 1669390400
transform 1 0 61152 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_537
timestamp 1669390400
transform 1 0 61488 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_80_601
timestamp 1669390400
transform 1 0 68656 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_80_665
timestamp 1669390400
transform 1 0 75824 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_80_681
timestamp 1669390400
transform 1 0 77616 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_80_685
timestamp 1669390400
transform 1 0 78064 0 1 65856
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_80_687
timestamp 1669390400
transform 1 0 78288 0 1 65856
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_2
timestamp 1669390400
transform 1 0 1568 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_66
timestamp 1669390400
transform 1 0 8736 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_130
timestamp 1669390400
transform 1 0 15904 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_194
timestamp 1669390400
transform 1 0 23072 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_258
timestamp 1669390400
transform 1 0 30240 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_81_322
timestamp 1669390400
transform 1 0 37408 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_81_354
timestamp 1669390400
transform 1 0 40992 0 -1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_356
timestamp 1669390400
transform 1 0 41216 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_359
timestamp 1669390400
transform 1 0 41552 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_423
timestamp 1669390400
transform 1 0 48720 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_487
timestamp 1669390400
transform 1 0 55888 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_551
timestamp 1669390400
transform 1 0 63056 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_81_615
timestamp 1669390400
transform 1 0 70224 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_81_679
timestamp 1669390400
transform 1 0 77392 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_81_687
timestamp 1669390400
transform 1 0 78288 0 -1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_2
timestamp 1669390400
transform 1 0 1568 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_66
timestamp 1669390400
transform 1 0 8736 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_82_130
timestamp 1669390400
transform 1 0 15904 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_82_162
timestamp 1669390400
transform 1 0 19488 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_180
timestamp 1669390400
transform 1 0 21504 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_244
timestamp 1669390400
transform 1 0 28672 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_308
timestamp 1669390400
transform 1 0 35840 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_372
timestamp 1669390400
transform 1 0 43008 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_436
timestamp 1669390400
transform 1 0 50176 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_82_500
timestamp 1669390400
transform 1 0 57344 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_532
timestamp 1669390400
transform 1 0 60928 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_534
timestamp 1669390400
transform 1 0 61152 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_537
timestamp 1669390400
transform 1 0 61488 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_82_601
timestamp 1669390400
transform 1 0 68656 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_82_665
timestamp 1669390400
transform 1 0 75824 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_82_681
timestamp 1669390400
transform 1 0 77616 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_82_685
timestamp 1669390400
transform 1 0 78064 0 1 67424
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_82_687
timestamp 1669390400
transform 1 0 78288 0 1 67424
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_2
timestamp 1669390400
transform 1 0 1568 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_66
timestamp 1669390400
transform 1 0 8736 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_130
timestamp 1669390400
transform 1 0 15904 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_194
timestamp 1669390400
transform 1 0 23072 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_258
timestamp 1669390400
transform 1 0 30240 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_83_322
timestamp 1669390400
transform 1 0 37408 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_83_354
timestamp 1669390400
transform 1 0 40992 0 -1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_356
timestamp 1669390400
transform 1 0 41216 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_359
timestamp 1669390400
transform 1 0 41552 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_423
timestamp 1669390400
transform 1 0 48720 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_487
timestamp 1669390400
transform 1 0 55888 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_551
timestamp 1669390400
transform 1 0 63056 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_83_615
timestamp 1669390400
transform 1 0 70224 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_83_679
timestamp 1669390400
transform 1 0 77392 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_83_687
timestamp 1669390400
transform 1 0 78288 0 -1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_2
timestamp 1669390400
transform 1 0 1568 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_66
timestamp 1669390400
transform 1 0 8736 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_84_130
timestamp 1669390400
transform 1 0 15904 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_84_162
timestamp 1669390400
transform 1 0 19488 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_180
timestamp 1669390400
transform 1 0 21504 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_244
timestamp 1669390400
transform 1 0 28672 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_84_308
timestamp 1669390400
transform 1 0 35840 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_324
timestamp 1669390400
transform 1 0 37632 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_328
timestamp 1669390400
transform 1 0 38080 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_330
timestamp 1669390400
transform 1 0 38304 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_333
timestamp 1669390400
transform 1 0 38640 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_337
timestamp 1669390400
transform 1 0 39088 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_343
timestamp 1669390400
transform 1 0 39760 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_84_347
timestamp 1669390400
transform 1 0 40208 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_84_363
timestamp 1669390400
transform 1 0 42000 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_371
timestamp 1669390400
transform 1 0 42896 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_84_375
timestamp 1669390400
transform 1 0 43344 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_383
timestamp 1669390400
transform 1 0 44240 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_386
timestamp 1669390400
transform 1 0 44576 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_390
timestamp 1669390400
transform 1 0 45024 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_84_454
timestamp 1669390400
transform 1 0 52192 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_470
timestamp 1669390400
transform 1 0 53984 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_474
timestamp 1669390400
transform 1 0 54432 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_84_477
timestamp 1669390400
transform 1 0 54768 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_84_509
timestamp 1669390400
transform 1 0 58352 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_84_525
timestamp 1669390400
transform 1 0 60144 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_533
timestamp 1669390400
transform 1 0 61040 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_537
timestamp 1669390400
transform 1 0 61488 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_84_601
timestamp 1669390400
transform 1 0 68656 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_84_665
timestamp 1669390400
transform 1 0 75824 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_84_681
timestamp 1669390400
transform 1 0 77616 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_84_685
timestamp 1669390400
transform 1 0 78064 0 1 68992
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_84_687
timestamp 1669390400
transform 1 0 78288 0 1 68992
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_2
timestamp 1669390400
transform 1 0 1568 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_66
timestamp 1669390400
transform 1 0 8736 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_130
timestamp 1669390400
transform 1 0 15904 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_194
timestamp 1669390400
transform 1 0 23072 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_85_258
timestamp 1669390400
transform 1 0 30240 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_85_290
timestamp 1669390400
transform 1 0 33824 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_85_306
timestamp 1669390400
transform 1 0 35616 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_314
timestamp 1669390400
transform 1 0 36512 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_318
timestamp 1669390400
transform 1 0 36960 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_321
timestamp 1669390400
transform 1 0 37296 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_325
timestamp 1669390400
transform 1 0 37744 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_329
timestamp 1669390400
transform 1 0 38192 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_333
timestamp 1669390400
transform 1 0 38640 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_337
timestamp 1669390400
transform 1 0 39088 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_343
timestamp 1669390400
transform 1 0 39760 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_345
timestamp 1669390400
transform 1 0 39984 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_351
timestamp 1669390400
transform 1 0 40656 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_355
timestamp 1669390400
transform 1 0 41104 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_85_359
timestamp 1669390400
transform 1 0 41552 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_367
timestamp 1669390400
transform 1 0 42448 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_377
timestamp 1669390400
transform 1 0 43568 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_381
timestamp 1669390400
transform 1 0 44016 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_385
timestamp 1669390400
transform 1 0 44464 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_389
timestamp 1669390400
transform 1 0 44912 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_393
timestamp 1669390400
transform 1 0 45360 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_397
timestamp 1669390400
transform 1 0 45808 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_401
timestamp 1669390400
transform 1 0 46256 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_405
timestamp 1669390400
transform 1 0 46704 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_407
timestamp 1669390400
transform 1 0 46928 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_85_410
timestamp 1669390400
transform 1 0 47264 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_426
timestamp 1669390400
transform 1 0 49056 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_430
timestamp 1669390400
transform 1 0 49504 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_433
timestamp 1669390400
transform 1 0 49840 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_437
timestamp 1669390400
transform 1 0 50288 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_441
timestamp 1669390400
transform 1 0 50736 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_445
timestamp 1669390400
transform 1 0 51184 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_447
timestamp 1669390400
transform 1 0 51408 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_450
timestamp 1669390400
transform 1 0 51744 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_454
timestamp 1669390400
transform 1 0 52192 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_458
timestamp 1669390400
transform 1 0 52640 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_462
timestamp 1669390400
transform 1 0 53088 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_466
timestamp 1669390400
transform 1 0 53536 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_470
timestamp 1669390400
transform 1 0 53984 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_473
timestamp 1669390400
transform 1 0 54320 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_477
timestamp 1669390400
transform 1 0 54768 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_483
timestamp 1669390400
transform 1 0 55440 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_489
timestamp 1669390400
transform 1 0 56112 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_493
timestamp 1669390400
transform 1 0 56560 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_497
timestamp 1669390400
transform 1 0 57008 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_85_561
timestamp 1669390400
transform 1 0 64176 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_85_625
timestamp 1669390400
transform 1 0 71344 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_85_657
timestamp 1669390400
transform 1 0 74928 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_85_673
timestamp 1669390400
transform 1 0 76720 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_85_681
timestamp 1669390400
transform 1 0 77616 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_85_685
timestamp 1669390400
transform 1 0 78064 0 -1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_85_687
timestamp 1669390400
transform 1 0 78288 0 -1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_2
timestamp 1669390400
transform 1 0 1568 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_66
timestamp 1669390400
transform 1 0 8736 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_86_130
timestamp 1669390400
transform 1 0 15904 0 1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_86_162
timestamp 1669390400
transform 1 0 19488 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_180
timestamp 1669390400
transform 1 0 21504 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_86_244
timestamp 1669390400
transform 1 0 28672 0 1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_86_276
timestamp 1669390400
transform 1 0 32256 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_86_292
timestamp 1669390400
transform 1 0 34048 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_300
timestamp 1669390400
transform 1 0 34944 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_303
timestamp 1669390400
transform 1 0 35280 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_307
timestamp 1669390400
transform 1 0 35728 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_311
timestamp 1669390400
transform 1 0 36176 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_315
timestamp 1669390400
transform 1 0 36624 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_319
timestamp 1669390400
transform 1 0 37072 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_322
timestamp 1669390400
transform 1 0 37408 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_326
timestamp 1669390400
transform 1 0 37856 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_330
timestamp 1669390400
transform 1 0 38304 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_338
timestamp 1669390400
transform 1 0 39200 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_347
timestamp 1669390400
transform 1 0 40208 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_362
timestamp 1669390400
transform 1 0 41888 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_366
timestamp 1669390400
transform 1 0 42336 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_368
timestamp 1669390400
transform 1 0 42560 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_393
timestamp 1669390400
transform 1 0 45360 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_397
timestamp 1669390400
transform 1 0 45808 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_401
timestamp 1669390400
transform 1 0 46256 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_405
timestamp 1669390400
transform 1 0 46704 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_409
timestamp 1669390400
transform 1 0 47152 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_413
timestamp 1669390400
transform 1 0 47600 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_417
timestamp 1669390400
transform 1 0 48048 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_421
timestamp 1669390400
transform 1 0 48496 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_425
timestamp 1669390400
transform 1 0 48944 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_429
timestamp 1669390400
transform 1 0 49392 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_433
timestamp 1669390400
transform 1 0 49840 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_439
timestamp 1669390400
transform 1 0 50512 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_443
timestamp 1669390400
transform 1 0 50960 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_447
timestamp 1669390400
transform 1 0 51408 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_457
timestamp 1669390400
transform 1 0 52528 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_461
timestamp 1669390400
transform 1 0 52976 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_465
timestamp 1669390400
transform 1 0 53424 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_469
timestamp 1669390400
transform 1 0 53872 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_472
timestamp 1669390400
transform 1 0 54208 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_476
timestamp 1669390400
transform 1 0 54656 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_480
timestamp 1669390400
transform 1 0 55104 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_484
timestamp 1669390400
transform 1 0 55552 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_494
timestamp 1669390400
transform 1 0 56672 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_502
timestamp 1669390400
transform 1 0 57568 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_86_506
timestamp 1669390400
transform 1 0 58016 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_86_522
timestamp 1669390400
transform 1 0 59808 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_530
timestamp 1669390400
transform 1 0 60704 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_534
timestamp 1669390400
transform 1 0 61152 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_537
timestamp 1669390400
transform 1 0 61488 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_86_601
timestamp 1669390400
transform 1 0 68656 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_86_665
timestamp 1669390400
transform 1 0 75824 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_86_681
timestamp 1669390400
transform 1 0 77616 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_86_685
timestamp 1669390400
transform 1 0 78064 0 1 70560
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_86_687
timestamp 1669390400
transform 1 0 78288 0 1 70560
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_2
timestamp 1669390400
transform 1 0 1568 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_66
timestamp 1669390400
transform 1 0 8736 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_130
timestamp 1669390400
transform 1 0 15904 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_194
timestamp 1669390400
transform 1 0 23072 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_87_258
timestamp 1669390400
transform 1 0 30240 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_292
timestamp 1669390400
transform 1 0 34048 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_296
timestamp 1669390400
transform 1 0 34496 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_302
timestamp 1669390400
transform 1 0 35168 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_306
timestamp 1669390400
transform 1 0 35616 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_310
timestamp 1669390400
transform 1 0 36064 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_314
timestamp 1669390400
transform 1 0 36512 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_320
timestamp 1669390400
transform 1 0 37184 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_327
timestamp 1669390400
transform 1 0 37968 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_352
timestamp 1669390400
transform 1 0 40768 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_356
timestamp 1669390400
transform 1 0 41216 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_359
timestamp 1669390400
transform 1 0 41552 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_383
timestamp 1669390400
transform 1 0 44240 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_393
timestamp 1669390400
transform 1 0 45360 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_399
timestamp 1669390400
transform 1 0 46032 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_403
timestamp 1669390400
transform 1 0 46480 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_407
timestamp 1669390400
transform 1 0 46928 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_411
timestamp 1669390400
transform 1 0 47376 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_415
timestamp 1669390400
transform 1 0 47824 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_419
timestamp 1669390400
transform 1 0 48272 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_423
timestamp 1669390400
transform 1 0 48720 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_427
timestamp 1669390400
transform 1 0 49168 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_452
timestamp 1669390400
transform 1 0 51968 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_458
timestamp 1669390400
transform 1 0 52640 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_472
timestamp 1669390400
transform 1 0 54208 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_476
timestamp 1669390400
transform 1 0 54656 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_87_478
timestamp 1669390400
transform 1 0 54880 0 -1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_485
timestamp 1669390400
transform 1 0 55664 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_510
timestamp 1669390400
transform 1 0 58464 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_514
timestamp 1669390400
transform 1 0 58912 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_518
timestamp 1669390400
transform 1 0 59360 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_522
timestamp 1669390400
transform 1 0 59808 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_87_586
timestamp 1669390400
transform 1 0 66976 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_87_650
timestamp 1669390400
transform 1 0 74144 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_87_682
timestamp 1669390400
transform 1 0 77728 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_87_686
timestamp 1669390400
transform 1 0 78176 0 -1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_2
timestamp 1669390400
transform 1 0 1568 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_66
timestamp 1669390400
transform 1 0 8736 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_88_130
timestamp 1669390400
transform 1 0 15904 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_88_162
timestamp 1669390400
transform 1 0 19488 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_180
timestamp 1669390400
transform 1 0 21504 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_88_244
timestamp 1669390400
transform 1 0 28672 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_88_260
timestamp 1669390400
transform 1 0 30464 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_268
timestamp 1669390400
transform 1 0 31360 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_274
timestamp 1669390400
transform 1 0 32032 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_278
timestamp 1669390400
transform 1 0 32480 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_282
timestamp 1669390400
transform 1 0 32928 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_286
timestamp 1669390400
transform 1 0 33376 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_290
timestamp 1669390400
transform 1 0 33824 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_294
timestamp 1669390400
transform 1 0 34272 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_300
timestamp 1669390400
transform 1 0 34944 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_306
timestamp 1669390400
transform 1 0 35616 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_310
timestamp 1669390400
transform 1 0 36064 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_315
timestamp 1669390400
transform 1 0 36624 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_329
timestamp 1669390400
transform 1 0 38192 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_333
timestamp 1669390400
transform 1 0 38640 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_358
timestamp 1669390400
transform 1 0 41440 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_362
timestamp 1669390400
transform 1 0 41888 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_376
timestamp 1669390400
transform 1 0 43456 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_384
timestamp 1669390400
transform 1 0 44352 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_398
timestamp 1669390400
transform 1 0 45920 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_405
timestamp 1669390400
transform 1 0 46704 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_411
timestamp 1669390400
transform 1 0 47376 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_415
timestamp 1669390400
transform 1 0 47824 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_421
timestamp 1669390400
transform 1 0 48496 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_423
timestamp 1669390400
transform 1 0 48720 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_428
timestamp 1669390400
transform 1 0 49280 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_438
timestamp 1669390400
transform 1 0 50400 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_444
timestamp 1669390400
transform 1 0 51072 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_446
timestamp 1669390400
transform 1 0 51296 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_470
timestamp 1669390400
transform 1 0 53984 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_480
timestamp 1669390400
transform 1 0 55104 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_487
timestamp 1669390400
transform 1 0 55888 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_489
timestamp 1669390400
transform 1 0 56112 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_513
timestamp 1669390400
transform 1 0 58800 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_519
timestamp 1669390400
transform 1 0 59472 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_523
timestamp 1669390400
transform 1 0 59920 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_527
timestamp 1669390400
transform 1 0 60368 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_531
timestamp 1669390400
transform 1 0 60816 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_537
timestamp 1669390400
transform 1 0 61488 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_88_601
timestamp 1669390400
transform 1 0 68656 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_88_665
timestamp 1669390400
transform 1 0 75824 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_88_681
timestamp 1669390400
transform 1 0 77616 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_88_685
timestamp 1669390400
transform 1 0 78064 0 1 72128
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_88_687
timestamp 1669390400
transform 1 0 78288 0 1 72128
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_2
timestamp 1669390400
transform 1 0 1568 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_66
timestamp 1669390400
transform 1 0 8736 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_130
timestamp 1669390400
transform 1 0 15904 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_194
timestamp 1669390400
transform 1 0 23072 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_258
timestamp 1669390400
transform 1 0 30240 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_261
timestamp 1669390400
transform 1 0 30576 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_265
timestamp 1669390400
transform 1 0 31024 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_271
timestamp 1669390400
transform 1 0 31696 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_273
timestamp 1669390400
transform 1 0 31920 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_276
timestamp 1669390400
transform 1 0 32256 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_282
timestamp 1669390400
transform 1 0 32928 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_290
timestamp 1669390400
transform 1 0 33824 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_298
timestamp 1669390400
transform 1 0 34720 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_306
timestamp 1669390400
transform 1 0 35616 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_313
timestamp 1669390400
transform 1 0 36400 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_320
timestamp 1669390400
transform 1 0 37184 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_328
timestamp 1669390400
transform 1 0 38080 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_338
timestamp 1669390400
transform 1 0 39200 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_346
timestamp 1669390400
transform 1 0 40096 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_356
timestamp 1669390400
transform 1 0 41216 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_359
timestamp 1669390400
transform 1 0 41552 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_362
timestamp 1669390400
transform 1 0 41888 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_364
timestamp 1669390400
transform 1 0 42112 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_375
timestamp 1669390400
transform 1 0 43344 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_379
timestamp 1669390400
transform 1 0 43792 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_391
timestamp 1669390400
transform 1 0 45136 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_405
timestamp 1669390400
transform 1 0 46704 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_412
timestamp 1669390400
transform 1 0 47488 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_418
timestamp 1669390400
transform 1 0 48160 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_424
timestamp 1669390400
transform 1 0 48832 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_438
timestamp 1669390400
transform 1 0 50400 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_446
timestamp 1669390400
transform 1 0 51296 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_89_448
timestamp 1669390400
transform 1 0 51520 0 -1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_462
timestamp 1669390400
transform 1 0 53088 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_472
timestamp 1669390400
transform 1 0 54208 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_480
timestamp 1669390400
transform 1 0 55104 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_484
timestamp 1669390400
transform 1 0 55552 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_89_494
timestamp 1669390400
transform 1 0 56672 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_510
timestamp 1669390400
transform 1 0 58464 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_524
timestamp 1669390400
transform 1 0 60032 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_530
timestamp 1669390400
transform 1 0 60704 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_534
timestamp 1669390400
transform 1 0 61152 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_538
timestamp 1669390400
transform 1 0 61600 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_542
timestamp 1669390400
transform 1 0 62048 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_89_606
timestamp 1669390400
transform 1 0 69216 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_89_670
timestamp 1669390400
transform 1 0 76384 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_89_686
timestamp 1669390400
transform 1 0 78176 0 -1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_2
timestamp 1669390400
transform 1 0 1568 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_66
timestamp 1669390400
transform 1 0 8736 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_90_130
timestamp 1669390400
transform 1 0 15904 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_90_162
timestamp 1669390400
transform 1 0 19488 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_180
timestamp 1669390400
transform 1 0 21504 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_244
timestamp 1669390400
transform 1 0 28672 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_247
timestamp 1669390400
transform 1 0 29008 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_251
timestamp 1669390400
transform 1 0 29456 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_255
timestamp 1669390400
transform 1 0 29904 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_263
timestamp 1669390400
transform 1 0 30800 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_271
timestamp 1669390400
transform 1 0 31696 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_279
timestamp 1669390400
transform 1 0 32592 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_281
timestamp 1669390400
transform 1 0 32816 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_288
timestamp 1669390400
transform 1 0 33600 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_298
timestamp 1669390400
transform 1 0 34720 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_308
timestamp 1669390400
transform 1 0 35840 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_325
timestamp 1669390400
transform 1 0 37744 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_331
timestamp 1669390400
transform 1 0 38416 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_341
timestamp 1669390400
transform 1 0 39536 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_345
timestamp 1669390400
transform 1 0 39984 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_355
timestamp 1669390400
transform 1 0 41104 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_376
timestamp 1669390400
transform 1 0 43456 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_386
timestamp 1669390400
transform 1 0 44576 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_390
timestamp 1669390400
transform 1 0 45024 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_392
timestamp 1669390400
transform 1 0 45248 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_401
timestamp 1669390400
transform 1 0 46256 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_407
timestamp 1669390400
transform 1 0 46928 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_413
timestamp 1669390400
transform 1 0 47600 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_417
timestamp 1669390400
transform 1 0 48048 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_419
timestamp 1669390400
transform 1 0 48272 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_425
timestamp 1669390400
transform 1 0 48944 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_437
timestamp 1669390400
transform 1 0 50288 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_448
timestamp 1669390400
transform 1 0 51520 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_455
timestamp 1669390400
transform 1 0 52304 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_474
timestamp 1669390400
transform 1 0 54432 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_481
timestamp 1669390400
transform 1 0 55216 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_483
timestamp 1669390400
transform 1 0 55440 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_489
timestamp 1669390400
transform 1 0 56112 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_493
timestamp 1669390400
transform 1 0 56560 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_500
timestamp 1669390400
transform 1 0 57344 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_507
timestamp 1669390400
transform 1 0 58128 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_519
timestamp 1669390400
transform 1 0 59472 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_525
timestamp 1669390400
transform 1 0 60144 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_90_531
timestamp 1669390400
transform 1 0 60816 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_537
timestamp 1669390400
transform 1 0 61488 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_540
timestamp 1669390400
transform 1 0 61824 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_544
timestamp 1669390400
transform 1 0 62272 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_548
timestamp 1669390400
transform 1 0 62720 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_90_552
timestamp 1669390400
transform 1 0 63168 0 1 73696
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_556
timestamp 1669390400
transform 1 0 63616 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_90_620
timestamp 1669390400
transform 1 0 70784 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_684
timestamp 1669390400
transform 1 0 77952 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_90_687
timestamp 1669390400
transform 1 0 78288 0 1 73696
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_2
timestamp 1669390400
transform 1 0 1568 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_66
timestamp 1669390400
transform 1 0 8736 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_91_130
timestamp 1669390400
transform 1 0 15904 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_91_194
timestamp 1669390400
transform 1 0 23072 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_91_226
timestamp 1669390400
transform 1 0 26656 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_246
timestamp 1669390400
transform 1 0 28896 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_252
timestamp 1669390400
transform 1 0 29568 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_260
timestamp 1669390400
transform 1 0 30464 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_270
timestamp 1669390400
transform 1 0 31584 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_272
timestamp 1669390400
transform 1 0 31808 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_281
timestamp 1669390400
transform 1 0 32816 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_291
timestamp 1669390400
transform 1 0 33936 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_299
timestamp 1669390400
transform 1 0 34832 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_309
timestamp 1669390400
transform 1 0 35952 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_326
timestamp 1669390400
transform 1 0 37856 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_338
timestamp 1669390400
transform 1 0 39200 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_348
timestamp 1669390400
transform 1 0 40320 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_356
timestamp 1669390400
transform 1 0 41216 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_359
timestamp 1669390400
transform 1 0 41552 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_362
timestamp 1669390400
transform 1 0 41888 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_364
timestamp 1669390400
transform 1 0 42112 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_375
timestamp 1669390400
transform 1 0 43344 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_387
timestamp 1669390400
transform 1 0 44688 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_391
timestamp 1669390400
transform 1 0 45136 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_393
timestamp 1669390400
transform 1 0 45360 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_404
timestamp 1669390400
transform 1 0 46592 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_411
timestamp 1669390400
transform 1 0 47376 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_415
timestamp 1669390400
transform 1 0 47824 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_431
timestamp 1669390400
transform 1 0 49616 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_439
timestamp 1669390400
transform 1 0 50512 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_441
timestamp 1669390400
transform 1 0 50736 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_454
timestamp 1669390400
transform 1 0 52192 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_456
timestamp 1669390400
transform 1 0 52416 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_463
timestamp 1669390400
transform 1 0 53200 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_475
timestamp 1669390400
transform 1 0 54544 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_487
timestamp 1669390400
transform 1 0 55888 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_506
timestamp 1669390400
transform 1 0 58016 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_510
timestamp 1669390400
transform 1 0 58464 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_522
timestamp 1669390400
transform 1 0 59808 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_528
timestamp 1669390400
transform 1 0 60480 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_534
timestamp 1669390400
transform 1 0 61152 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_540
timestamp 1669390400
transform 1 0 61824 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_546
timestamp 1669390400
transform 1 0 62496 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_552
timestamp 1669390400
transform 1 0 63168 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_556
timestamp 1669390400
transform 1 0 63616 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_91_560
timestamp 1669390400
transform 1 0 64064 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_576
timestamp 1669390400
transform 1 0 65856 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_580
timestamp 1669390400
transform 1 0 66304 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_582
timestamp 1669390400
transform 1 0 66528 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_585
timestamp 1669390400
transform 1 0 66864 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_589
timestamp 1669390400
transform 1 0 67312 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_91_595
timestamp 1669390400
transform 1 0 67984 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_91_611
timestamp 1669390400
transform 1 0 69776 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_91_621
timestamp 1669390400
transform 1 0 70896 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_91_639
timestamp 1669390400
transform 1 0 72912 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_647
timestamp 1669390400
transform 1 0 73808 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_91_655
timestamp 1669390400
transform 1 0 74704 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_667
timestamp 1669390400
transform 1 0 76048 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_91_673
timestamp 1669390400
transform 1 0 76720 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_677
timestamp 1669390400
transform 1 0 77168 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_91_681
timestamp 1669390400
transform 1 0 77616 0 -1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_91_687
timestamp 1669390400
transform 1 0 78288 0 -1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_2
timestamp 1669390400
transform 1 0 1568 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_5
timestamp 1669390400
transform 1 0 1904 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_13
timestamp 1669390400
transform 1 0 2800 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_19
timestamp 1669390400
transform 1 0 3472 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_27
timestamp 1669390400
transform 1 0 4368 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_31
timestamp 1669390400
transform 1 0 4816 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_92_37
timestamp 1669390400
transform 1 0 5488 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_101
timestamp 1669390400
transform 1 0 12656 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_109
timestamp 1669390400
transform 1 0 13552 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_113
timestamp 1669390400
transform 1 0 14000 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_121
timestamp 1669390400
transform 1 0 14896 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_127
timestamp 1669390400
transform 1 0 15568 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_131
timestamp 1669390400
transform 1 0 16016 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_139
timestamp 1669390400
transform 1 0 16912 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_145
timestamp 1669390400
transform 1 0 17584 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_149
timestamp 1669390400
transform 1 0 18032 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_157
timestamp 1669390400
transform 1 0 18928 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_163
timestamp 1669390400
transform 1 0 19600 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_167
timestamp 1669390400
transform 1 0 20048 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_177
timestamp 1669390400
transform 1 0 21168 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_180
timestamp 1669390400
transform 1 0 21504 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_185
timestamp 1669390400
transform 1 0 22064 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_193
timestamp 1669390400
transform 1 0 22960 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_199
timestamp 1669390400
transform 1 0 23632 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_203
timestamp 1669390400
transform 1 0 24080 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_211
timestamp 1669390400
transform 1 0 24976 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_92_217
timestamp 1669390400
transform 1 0 25648 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_225
timestamp 1669390400
transform 1 0 26544 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_229
timestamp 1669390400
transform 1 0 26992 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_235
timestamp 1669390400
transform 1 0 27664 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_245
timestamp 1669390400
transform 1 0 28784 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_253
timestamp 1669390400
transform 1 0 29680 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_263
timestamp 1669390400
transform 1 0 30800 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_273
timestamp 1669390400
transform 1 0 31920 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_281
timestamp 1669390400
transform 1 0 32816 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_291
timestamp 1669390400
transform 1 0 33936 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_297
timestamp 1669390400
transform 1 0 34608 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_307
timestamp 1669390400
transform 1 0 35728 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_309
timestamp 1669390400
transform 1 0 35952 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_319
timestamp 1669390400
transform 1 0 37072 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_325
timestamp 1669390400
transform 1 0 37744 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_341
timestamp 1669390400
transform 1 0 39536 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_353
timestamp 1669390400
transform 1 0 40880 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_362
timestamp 1669390400
transform 1 0 41888 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_373
timestamp 1669390400
transform 1 0 43120 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_384
timestamp 1669390400
transform 1 0 44352 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_392
timestamp 1669390400
transform 1 0 45248 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_400
timestamp 1669390400
transform 1 0 46144 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_408
timestamp 1669390400
transform 1 0 47040 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_416
timestamp 1669390400
transform 1 0 47936 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_422
timestamp 1669390400
transform 1 0 48608 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_434
timestamp 1669390400
transform 1 0 49952 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_446
timestamp 1669390400
transform 1 0 51296 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_456
timestamp 1669390400
transform 1 0 52416 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_464
timestamp 1669390400
transform 1 0 53312 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_476
timestamp 1669390400
transform 1 0 54656 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_486
timestamp 1669390400
transform 1 0 55776 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_494
timestamp 1669390400
transform 1 0 56672 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_502
timestamp 1669390400
transform 1 0 57568 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_510
timestamp 1669390400
transform 1 0 58464 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_518
timestamp 1669390400
transform 1 0 59360 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_525
timestamp 1669390400
transform 1 0 60144 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_531
timestamp 1669390400
transform 1 0 60816 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_537
timestamp 1669390400
transform 1 0 61488 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_542
timestamp 1669390400
transform 1 0 62048 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_548
timestamp 1669390400
transform 1 0 62720 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_554
timestamp 1669390400
transform 1 0 63392 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_560
timestamp 1669390400
transform 1 0 64064 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_566
timestamp 1669390400
transform 1 0 64736 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_568
timestamp 1669390400
transform 1 0 64960 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_571
timestamp 1669390400
transform 1 0 65296 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_577
timestamp 1669390400
transform 1 0 65968 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_583
timestamp 1669390400
transform 1 0 66640 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_610
timestamp 1669390400
transform 1 0 69664 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_616
timestamp 1669390400
transform 1 0 70336 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_622
timestamp 1669390400
transform 1 0 71008 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_626
timestamp 1669390400
transform 1 0 71456 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_631
timestamp 1669390400
transform 1 0 72016 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_637
timestamp 1669390400
transform 1 0 72688 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_645
timestamp 1669390400
transform 1 0 73584 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_92_651
timestamp 1669390400
transform 1 0 74256 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_655
timestamp 1669390400
transform 1 0 74704 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_92_681
timestamp 1669390400
transform 1 0 77616 0 1 75264
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_92_687
timestamp 1669390400
transform 1 0 78288 0 1 75264
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_2
timestamp 1669390400
transform 1 0 1568 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_19
timestamp 1669390400
transform 1 0 3472 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_35
timestamp 1669390400
transform 1 0 5264 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_43
timestamp 1669390400
transform 1 0 6160 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_47
timestamp 1669390400
transform 1 0 6608 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_55
timestamp 1669390400
transform 1 0 7504 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_93_61
timestamp 1669390400
transform 1 0 8176 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_73
timestamp 1669390400
transform 1 0 9520 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_93_79
timestamp 1669390400
transform 1 0 10192 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_91
timestamp 1669390400
transform 1 0 11536 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_107
timestamp 1669390400
transform 1 0 13328 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_125
timestamp 1669390400
transform 1 0 15344 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_143
timestamp 1669390400
transform 1 0 17360 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_161
timestamp 1669390400
transform 1 0 19376 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_177
timestamp 1669390400
transform 1 0 21168 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_180
timestamp 1669390400
transform 1 0 21504 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_182
timestamp 1669390400
transform 1 0 21728 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_197
timestamp 1669390400
transform 1 0 23408 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_215
timestamp 1669390400
transform 1 0 25424 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_233
timestamp 1669390400
transform 1 0 27440 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_251
timestamp 1669390400
transform 1 0 29456 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_269
timestamp 1669390400
transform 1 0 31472 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_287
timestamp 1669390400
transform 1 0 33488 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_305
timestamp 1669390400
transform 1 0 35504 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_323
timestamp 1669390400
transform 1 0 37520 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_331
timestamp 1669390400
transform 1 0 38416 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_349
timestamp 1669390400
transform 1 0 40432 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_355
timestamp 1669390400
transform 1 0 41104 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_358
timestamp 1669390400
transform 1 0 41440 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_375
timestamp 1669390400
transform 1 0 43344 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_383
timestamp 1669390400
transform 1 0 44240 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_391
timestamp 1669390400
transform 1 0 45136 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_399
timestamp 1669390400
transform 1 0 46032 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_403
timestamp 1669390400
transform 1 0 46480 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_430
timestamp 1669390400
transform 1 0 49504 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_439
timestamp 1669390400
transform 1 0 50512 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_466
timestamp 1669390400
transform 1 0 53536 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_474
timestamp 1669390400
transform 1 0 54432 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_476
timestamp 1669390400
transform 1 0 54656 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_493
timestamp 1669390400
transform 1 0 56560 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_511
timestamp 1669390400
transform 1 0 58576 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_519
timestamp 1669390400
transform 1 0 59472 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_525
timestamp 1669390400
transform 1 0 60144 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_531
timestamp 1669390400
transform 1 0 60816 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_533
timestamp 1669390400
transform 1 0 61040 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_536
timestamp 1669390400
transform 1 0 61376 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_543
timestamp 1669390400
transform 1 0 62160 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_547
timestamp 1669390400
transform 1 0 62608 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_574
timestamp 1669390400
transform 1 0 65632 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_601
timestamp 1669390400
transform 1 0 68656 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_609
timestamp 1669390400
transform 1 0 69552 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_615
timestamp 1669390400
transform 1 0 70224 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_619
timestamp 1669390400
transform 1 0 70672 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_93_646
timestamp 1669390400
transform 1 0 73696 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_93_650
timestamp 1669390400
transform 1 0 74144 0 -1 76832
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_652
timestamp 1669390400
transform 1 0 74368 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_93_687
timestamp 1669390400
transform 1 0 78288 0 -1 76832
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 78624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 78624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 78624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 78624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 78624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 78624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 78624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 78624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 78624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 78624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 78624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 78624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1669390400
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1669390400
transform -1 0 78624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1669390400
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1669390400
transform -1 0 78624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1669390400
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1669390400
transform -1 0 78624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1669390400
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1669390400
transform -1 0 78624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1669390400
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1669390400
transform -1 0 78624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1669390400
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1669390400
transform -1 0 78624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1669390400
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1669390400
transform -1 0 78624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1669390400
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1669390400
transform -1 0 78624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1669390400
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1669390400
transform -1 0 78624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1669390400
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1669390400
transform -1 0 78624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1669390400
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1669390400
transform -1 0 78624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1669390400
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1669390400
transform -1 0 78624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1669390400
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1669390400
transform -1 0 78624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1669390400
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1669390400
transform -1 0 78624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1669390400
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1669390400
transform -1 0 78624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1669390400
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1669390400
transform -1 0 78624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1669390400
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1669390400
transform -1 0 78624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1669390400
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1669390400
transform -1 0 78624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1669390400
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1669390400
transform -1 0 78624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1669390400
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1669390400
transform -1 0 78624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1669390400
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1669390400
transform -1 0 78624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1669390400
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1669390400
transform -1 0 78624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1669390400
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1669390400
transform -1 0 78624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1669390400
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1669390400
transform -1 0 78624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1669390400
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1669390400
transform -1 0 78624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1669390400
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1669390400
transform -1 0 78624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1669390400
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1669390400
transform -1 0 78624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1669390400
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1669390400
transform -1 0 78624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1669390400
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1669390400
transform -1 0 78624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1669390400
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1669390400
transform -1 0 78624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1669390400
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1669390400
transform -1 0 78624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1669390400
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1669390400
transform -1 0 78624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1669390400
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1669390400
transform -1 0 78624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1669390400
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1669390400
transform -1 0 78624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1669390400
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1669390400
transform -1 0 78624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1669390400
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1669390400
transform -1 0 78624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1669390400
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1669390400
transform -1 0 78624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1669390400
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1669390400
transform -1 0 78624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1669390400
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1669390400
transform -1 0 78624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1669390400
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1669390400
transform -1 0 78624 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1669390400
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1669390400
transform -1 0 78624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1669390400
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1669390400
transform -1 0 78624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1669390400
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1669390400
transform -1 0 78624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_110
timestamp 1669390400
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_111
timestamp 1669390400
transform -1 0 78624 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_112
timestamp 1669390400
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_113
timestamp 1669390400
transform -1 0 78624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_114
timestamp 1669390400
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_115
timestamp 1669390400
transform -1 0 78624 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_116
timestamp 1669390400
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_117
timestamp 1669390400
transform -1 0 78624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_118
timestamp 1669390400
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_119
timestamp 1669390400
transform -1 0 78624 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_120
timestamp 1669390400
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_121
timestamp 1669390400
transform -1 0 78624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_122
timestamp 1669390400
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_123
timestamp 1669390400
transform -1 0 78624 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_124
timestamp 1669390400
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_125
timestamp 1669390400
transform -1 0 78624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_126
timestamp 1669390400
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_127
timestamp 1669390400
transform -1 0 78624 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_128
timestamp 1669390400
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_129
timestamp 1669390400
transform -1 0 78624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_130
timestamp 1669390400
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_131
timestamp 1669390400
transform -1 0 78624 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_132
timestamp 1669390400
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_133
timestamp 1669390400
transform -1 0 78624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_134
timestamp 1669390400
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_135
timestamp 1669390400
transform -1 0 78624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_136
timestamp 1669390400
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_137
timestamp 1669390400
transform -1 0 78624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_138
timestamp 1669390400
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_139
timestamp 1669390400
transform -1 0 78624 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_140
timestamp 1669390400
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_141
timestamp 1669390400
transform -1 0 78624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_142
timestamp 1669390400
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_143
timestamp 1669390400
transform -1 0 78624 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_144
timestamp 1669390400
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_145
timestamp 1669390400
transform -1 0 78624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_146
timestamp 1669390400
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_147
timestamp 1669390400
transform -1 0 78624 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_148
timestamp 1669390400
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_149
timestamp 1669390400
transform -1 0 78624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_150
timestamp 1669390400
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_151
timestamp 1669390400
transform -1 0 78624 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_152
timestamp 1669390400
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_153
timestamp 1669390400
transform -1 0 78624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_154
timestamp 1669390400
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_155
timestamp 1669390400
transform -1 0 78624 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_156
timestamp 1669390400
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_157
timestamp 1669390400
transform -1 0 78624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_158
timestamp 1669390400
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_159
timestamp 1669390400
transform -1 0 78624 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_160
timestamp 1669390400
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_161
timestamp 1669390400
transform -1 0 78624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_162
timestamp 1669390400
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_163
timestamp 1669390400
transform -1 0 78624 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_164
timestamp 1669390400
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_165
timestamp 1669390400
transform -1 0 78624 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_166
timestamp 1669390400
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_167
timestamp 1669390400
transform -1 0 78624 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_168
timestamp 1669390400
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_169
timestamp 1669390400
transform -1 0 78624 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_170
timestamp 1669390400
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_171
timestamp 1669390400
transform -1 0 78624 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_172
timestamp 1669390400
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_173
timestamp 1669390400
transform -1 0 78624 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_174
timestamp 1669390400
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_175
timestamp 1669390400
transform -1 0 78624 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_176
timestamp 1669390400
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_177
timestamp 1669390400
transform -1 0 78624 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_178
timestamp 1669390400
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_179
timestamp 1669390400
transform -1 0 78624 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_180
timestamp 1669390400
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_181
timestamp 1669390400
transform -1 0 78624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_182
timestamp 1669390400
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_183
timestamp 1669390400
transform -1 0 78624 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_184
timestamp 1669390400
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_185
timestamp 1669390400
transform -1 0 78624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_186
timestamp 1669390400
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_187
timestamp 1669390400
transform -1 0 78624 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 21280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1669390400
transform 1 0 41216 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1669390400
transform 1 0 61152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1669390400
transform 1 0 41328 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1669390400
transform 1 0 21280 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1669390400
transform 1 0 61264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1669390400
transform 1 0 41328 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1669390400
transform 1 0 21280 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1669390400
transform 1 0 61264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1669390400
transform 1 0 41328 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1669390400
transform 1 0 21280 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1669390400
transform 1 0 61264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1669390400
transform 1 0 41328 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1669390400
transform 1 0 21280 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1669390400
transform 1 0 61264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1669390400
transform 1 0 41328 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1669390400
transform 1 0 21280 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1669390400
transform 1 0 61264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1669390400
transform 1 0 41328 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1669390400
transform 1 0 21280 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1669390400
transform 1 0 61264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1669390400
transform 1 0 41328 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1669390400
transform 1 0 21280 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1669390400
transform 1 0 61264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1669390400
transform 1 0 41328 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1669390400
transform 1 0 21280 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1669390400
transform 1 0 61264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1669390400
transform 1 0 41328 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1669390400
transform 1 0 21280 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1669390400
transform 1 0 61264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1669390400
transform 1 0 41328 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1669390400
transform 1 0 21280 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1669390400
transform 1 0 61264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1669390400
transform 1 0 41328 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1669390400
transform 1 0 21280 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1669390400
transform 1 0 61264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1669390400
transform 1 0 41328 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1669390400
transform 1 0 21280 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1669390400
transform 1 0 61264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1669390400
transform 1 0 41328 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1669390400
transform 1 0 21280 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1669390400
transform 1 0 61264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1669390400
transform 1 0 41328 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1669390400
transform 1 0 21280 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1669390400
transform 1 0 61264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1669390400
transform 1 0 41328 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1669390400
transform 1 0 21280 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1669390400
transform 1 0 61264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1669390400
transform 1 0 41328 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1669390400
transform 1 0 21280 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1669390400
transform 1 0 61264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1669390400
transform 1 0 41328 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1669390400
transform 1 0 21280 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1669390400
transform 1 0 61264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1669390400
transform 1 0 41328 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1669390400
transform 1 0 21280 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1669390400
transform 1 0 61264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1669390400
transform 1 0 41328 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1669390400
transform 1 0 21280 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1669390400
transform 1 0 61264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1669390400
transform 1 0 41328 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1669390400
transform 1 0 21280 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1669390400
transform 1 0 61264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1669390400
transform 1 0 41328 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1669390400
transform 1 0 21280 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1669390400
transform 1 0 61264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1669390400
transform 1 0 41328 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1669390400
transform 1 0 21280 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1669390400
transform 1 0 61264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1669390400
transform 1 0 41328 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1669390400
transform 1 0 21280 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1669390400
transform 1 0 61264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1669390400
transform 1 0 41328 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1669390400
transform 1 0 21280 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1669390400
transform 1 0 61264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1669390400
transform 1 0 41328 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1669390400
transform 1 0 21280 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1669390400
transform 1 0 61264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1669390400
transform 1 0 41328 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1669390400
transform 1 0 21280 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1669390400
transform 1 0 61264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1669390400
transform 1 0 41328 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1669390400
transform 1 0 21280 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1669390400
transform 1 0 61264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1669390400
transform 1 0 41328 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1669390400
transform 1 0 21280 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1669390400
transform 1 0 61264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1669390400
transform 1 0 41328 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1669390400
transform 1 0 21280 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1669390400
transform 1 0 61264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1669390400
transform 1 0 41328 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1669390400
transform 1 0 21280 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1669390400
transform 1 0 61264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1669390400
transform 1 0 41328 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1669390400
transform 1 0 21280 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1669390400
transform 1 0 61264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1669390400
transform 1 0 41328 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1669390400
transform 1 0 21280 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1669390400
transform 1 0 61264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1669390400
transform 1 0 41328 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1669390400
transform 1 0 21280 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1669390400
transform 1 0 61264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1669390400
transform 1 0 41328 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1669390400
transform 1 0 21280 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1669390400
transform 1 0 61264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1669390400
transform 1 0 41328 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1669390400
transform 1 0 21280 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1669390400
transform 1 0 61264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1669390400
transform 1 0 41328 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1669390400
transform 1 0 21280 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1669390400
transform 1 0 61264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1669390400
transform 1 0 41328 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1669390400
transform 1 0 21280 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1669390400
transform 1 0 61264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1669390400
transform 1 0 41328 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1669390400
transform 1 0 21280 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1669390400
transform 1 0 61264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1669390400
transform 1 0 41328 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1669390400
transform 1 0 21280 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1669390400
transform 1 0 61264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1669390400
transform 1 0 41328 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1669390400
transform 1 0 21280 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1669390400
transform 1 0 61264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1669390400
transform 1 0 41328 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1669390400
transform 1 0 21280 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1669390400
transform 1 0 61264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1669390400
transform 1 0 41328 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1669390400
transform 1 0 21280 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1669390400
transform 1 0 61264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1669390400
transform 1 0 41328 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1669390400
transform 1 0 21280 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1669390400
transform 1 0 61264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1669390400
transform 1 0 41328 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1669390400
transform 1 0 21280 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1669390400
transform 1 0 61264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1669390400
transform 1 0 41328 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1669390400
transform 1 0 21280 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1669390400
transform 1 0 61264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1669390400
transform 1 0 41328 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1669390400
transform 1 0 21280 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1669390400
transform 1 0 61264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1669390400
transform 1 0 21280 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1669390400
transform 1 0 41216 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1669390400
transform 1 0 61152 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _119_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 48608 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _120_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 46144 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _121_
timestamp 1669390400
transform 1 0 40544 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _122_
timestamp 1669390400
transform -1 0 47040 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _123_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 47376 0 -1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _124_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 45136 0 -1 73696
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _125_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 45920 0 1 72128
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _126_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 44352 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _127_
timestamp 1669390400
transform -1 0 48160 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _128_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 46592 0 -1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _129_
timestamp 1669390400
transform -1 0 46704 0 -1 73696
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _130_
timestamp 1669390400
transform -1 0 43456 0 1 72128
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _131_
timestamp 1669390400
transform -1 0 39760 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _132_
timestamp 1669390400
transform -1 0 39200 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _133_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 45360 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _134_
timestamp 1669390400
transform -1 0 40096 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _135_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 38304 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _136_
timestamp 1669390400
transform 1 0 37968 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _137_
timestamp 1669390400
transform -1 0 44240 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _138_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 40768 0 -1 72128
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _139_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 38864 0 1 72128
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _140_
timestamp 1669390400
transform -1 0 43568 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _141_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 41664 0 -1 72128
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1669390400
transform 1 0 46144 0 1 72128
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _143_
timestamp 1669390400
transform -1 0 47488 0 -1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _144_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 43344 0 -1 73696
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _145_
timestamp 1669390400
transform -1 0 41216 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _146_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 42224 0 -1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _147_
timestamp 1669390400
transform -1 0 60480 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _148_
timestamp 1669390400
transform -1 0 56672 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _149_
timestamp 1669390400
transform -1 0 53200 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _150_
timestamp 1669390400
transform -1 0 60144 0 1 75264
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _151_
timestamp 1669390400
transform -1 0 59360 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _152_
timestamp 1669390400
transform -1 0 55888 0 -1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _153_
timestamp 1669390400
transform -1 0 55216 0 1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _154_
timestamp 1669390400
transform -1 0 52192 0 -1 75264
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _155_
timestamp 1669390400
transform -1 0 51296 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _156_
timestamp 1669390400
transform -1 0 61824 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _157_
timestamp 1669390400
transform 1 0 58688 0 -1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _158_
timestamp 1669390400
transform -1 0 60032 0 -1 73696
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _159_
timestamp 1669390400
transform -1 0 54208 0 -1 72128
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _160_
timestamp 1669390400
transform -1 0 59472 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _161_
timestamp 1669390400
transform 1 0 54992 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _162_
timestamp 1669390400
transform 1 0 58576 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _163_
timestamp 1669390400
transform -1 0 57568 0 1 70560
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _164_
timestamp 1669390400
transform 1 0 55776 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _165_
timestamp 1669390400
transform -1 0 61152 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _166_
timestamp 1669390400
transform 1 0 56672 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _167_
timestamp 1669390400
transform 1 0 55888 0 -1 72128
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _168_
timestamp 1669390400
transform 1 0 56224 0 1 72128
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _169_
timestamp 1669390400
transform -1 0 55104 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _170_
timestamp 1669390400
transform -1 0 53984 0 1 72128
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _171_
timestamp 1669390400
transform 1 0 51520 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _172_
timestamp 1669390400
transform -1 0 51072 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _173_
timestamp 1669390400
transform 1 0 49280 0 -1 73696
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _174_
timestamp 1669390400
transform 1 0 49504 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _175_
timestamp 1669390400
transform -1 0 50288 0 1 73696
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _176_
timestamp 1669390400
transform 1 0 31024 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _177_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 50512 0 1 73696
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _178_
timestamp 1669390400
transform 1 0 42112 0 1 75264
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _179_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 43344 0 1 75264
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _180_
timestamp 1669390400
transform -1 0 35168 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _181_
timestamp 1669390400
transform -1 0 35616 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _182_
timestamp 1669390400
transform 1 0 35840 0 -1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _183_
timestamp 1669390400
transform 1 0 44576 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _184_
timestamp 1669390400
transform -1 0 46032 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _185_
timestamp 1669390400
transform -1 0 40320 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _186_
timestamp 1669390400
transform -1 0 40880 0 1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _187_
timestamp 1669390400
transform -1 0 55888 0 1 72128
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _188_
timestamp 1669390400
transform -1 0 53312 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _189_
timestamp 1669390400
transform -1 0 57568 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _190_
timestamp 1669390400
transform 1 0 54880 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _191_
timestamp 1669390400
transform -1 0 54656 0 1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _192_
timestamp 1669390400
transform 1 0 29792 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _193_
timestamp 1669390400
transform -1 0 30800 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _194_
timestamp 1669390400
transform -1 0 30800 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _195_
timestamp 1669390400
transform 1 0 31024 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _196_
timestamp 1669390400
transform 1 0 31920 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _197_
timestamp 1669390400
transform -1 0 29680 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _198_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 31584 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _199_
timestamp 1669390400
transform -1 0 38192 0 1 72128
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _200_
timestamp 1669390400
transform 1 0 38640 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _201_
timestamp 1669390400
transform -1 0 37968 0 -1 72128
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _202_
timestamp 1669390400
transform -1 0 37184 0 -1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _203_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 38416 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _204_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 36064 0 1 73696
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _205_
timestamp 1669390400
transform -1 0 58464 0 -1 73696
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _206_
timestamp 1669390400
transform 1 0 55776 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _207_
timestamp 1669390400
transform 1 0 55552 0 1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _208_
timestamp 1669390400
transform -1 0 58128 0 1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _209_
timestamp 1669390400
transform -1 0 58464 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _210_
timestamp 1669390400
transform 1 0 56336 0 -1 75264
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _211_
timestamp 1669390400
transform 1 0 31920 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _212_
timestamp 1669390400
transform 1 0 32928 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _213_
timestamp 1669390400
transform -1 0 33936 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _214_
timestamp 1669390400
transform 1 0 32144 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _215_
timestamp 1669390400
transform -1 0 33824 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _216_
timestamp 1669390400
transform 1 0 33040 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _217_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 40432 0 1 70560
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _218_
timestamp 1669390400
transform 1 0 37408 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _219_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 43568 0 -1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _220_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 44576 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _221_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 41552 0 1 73696
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _222_
timestamp 1669390400
transform 1 0 51632 0 -1 73696
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _223_
timestamp 1669390400
transform -1 0 55104 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _224_
timestamp 1669390400
transform 1 0 53424 0 -1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _225_
timestamp 1669390400
transform 1 0 53312 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _226_
timestamp 1669390400
transform 1 0 52528 0 1 73696
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _227_
timestamp 1669390400
transform 1 0 34048 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _228_
timestamp 1669390400
transform -1 0 35952 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _229_
timestamp 1669390400
transform 1 0 34832 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _230_
timestamp 1669390400
transform 1 0 44464 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _231_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 45360 0 1 70560
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _232_
timestamp 1669390400
transform 1 0 39648 0 1 70560
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _233_
timestamp 1669390400
transform 1 0 40208 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _234_
timestamp 1669390400
transform -1 0 40656 0 -1 70560
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _235_
timestamp 1669390400
transform 1 0 36176 0 -1 75264
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _236_
timestamp 1669390400
transform 1 0 51632 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _237_
timestamp 1669390400
transform -1 0 51968 0 -1 72128
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _238_
timestamp 1669390400
transform -1 0 52304 0 1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _239_
timestamp 1669390400
transform -1 0 51296 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _240_
timestamp 1669390400
transform -1 0 48944 0 1 73696
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _241_
timestamp 1669390400
transform 1 0 47936 0 -1 75264
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _242_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 50512 0 -1 76832
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _243_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 49952 0 1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _244_
timestamp 1669390400
transform -1 0 41888 0 1 75264
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _245_
timestamp 1669390400
transform -1 0 39200 0 -1 75264
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _246_
timestamp 1669390400
transform -1 0 37072 0 1 75264
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _247_
timestamp 1669390400
transform -1 0 34720 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _248_
timestamp 1669390400
transform -1 0 28784 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _249_
timestamp 1669390400
transform 1 0 29120 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _250_
timestamp 1669390400
transform -1 0 35840 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _251_
timestamp 1669390400
transform 1 0 34160 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _252_
timestamp 1669390400
transform 1 0 35168 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input1 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1680 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input2
timestamp 1669390400
transform 1 0 38640 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input3
timestamp 1669390400
transform -1 0 43344 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1669390400
transform -1 0 45136 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input5
timestamp 1669390400
transform 1 0 47264 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input6 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 49504 0 -1 76832
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1669390400
transform -1 0 50512 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input8
timestamp 1669390400
transform -1 0 53536 0 -1 76832
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input9
timestamp 1669390400
transform -1 0 54432 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input10
timestamp 1669390400
transform 1 0 54768 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input11
timestamp 1669390400
transform -1 0 58576 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1669390400
transform -1 0 59472 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input13
timestamp 1669390400
transform -1 0 62160 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input14
timestamp 1669390400
transform -1 0 65632 0 -1 76832
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input15
timestamp 1669390400
transform -1 0 68656 0 -1 76832
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input16
timestamp 1669390400
transform -1 0 69664 0 1 75264
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input17
timestamp 1669390400
transform -1 0 69552 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input18
timestamp 1669390400
transform -1 0 73696 0 -1 76832
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1669390400
transform -1 0 73584 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input20
timestamp 1669390400
transform -1 0 77616 0 1 75264
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyd_1  input21 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 78288 0 -1 76832
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_37 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 55440 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_38
timestamp 1669390400
transform -1 0 56112 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_39
timestamp 1669390400
transform -1 0 56784 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_40
timestamp 1669390400
transform -1 0 57456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_41
timestamp 1669390400
transform -1 0 58128 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_42
timestamp 1669390400
transform -1 0 58800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_43
timestamp 1669390400
transform -1 0 59472 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_44
timestamp 1669390400
transform -1 0 60144 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_45
timestamp 1669390400
transform -1 0 60816 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_46
timestamp 1669390400
transform -1 0 61936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_47
timestamp 1669390400
transform -1 0 62608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_48
timestamp 1669390400
transform -1 0 63280 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_49
timestamp 1669390400
transform -1 0 63952 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_50
timestamp 1669390400
transform -1 0 64624 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_51
timestamp 1669390400
transform -1 0 65296 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_52
timestamp 1669390400
transform -1 0 65968 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_53
timestamp 1669390400
transform -1 0 66640 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_54
timestamp 1669390400
transform -1 0 67312 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_55
timestamp 1669390400
transform -1 0 67984 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_56
timestamp 1669390400
transform -1 0 68656 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_57
timestamp 1669390400
transform -1 0 69328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_58
timestamp 1669390400
transform -1 0 70000 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_59
timestamp 1669390400
transform -1 0 70672 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_60
timestamp 1669390400
transform -1 0 71344 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_61
timestamp 1669390400
transform -1 0 72016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_62
timestamp 1669390400
transform -1 0 72688 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_63
timestamp 1669390400
transform -1 0 73360 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_64
timestamp 1669390400
transform -1 0 74032 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_65
timestamp 1669390400
transform -1 0 7280 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_66
timestamp 1669390400
transform -1 0 8624 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_67
timestamp 1669390400
transform -1 0 9520 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_68
timestamp 1669390400
transform -1 0 10416 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_69
timestamp 1669390400
transform -1 0 11088 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_70
timestamp 1669390400
transform 1 0 11312 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_71
timestamp 1669390400
transform 1 0 11984 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_72
timestamp 1669390400
transform 1 0 12656 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_73
timestamp 1669390400
transform 1 0 13328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_74
timestamp 1669390400
transform 1 0 14000 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_75
timestamp 1669390400
transform 1 0 14672 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_76
timestamp 1669390400
transform 1 0 15344 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_77
timestamp 1669390400
transform 1 0 16016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_78
timestamp 1669390400
transform 1 0 16688 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_79
timestamp 1669390400
transform 1 0 17360 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_80
timestamp 1669390400
transform 1 0 18032 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_81
timestamp 1669390400
transform 1 0 18704 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_82
timestamp 1669390400
transform 1 0 19376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_83
timestamp 1669390400
transform 1 0 20048 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_84
timestamp 1669390400
transform 1 0 20720 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_85
timestamp 1669390400
transform -1 0 22064 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_86
timestamp 1669390400
transform -1 0 22736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_87
timestamp 1669390400
transform -1 0 23408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_88
timestamp 1669390400
transform -1 0 24080 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_89
timestamp 1669390400
transform -1 0 24752 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_90
timestamp 1669390400
transform -1 0 25424 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_91
timestamp 1669390400
transform -1 0 26096 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_92
timestamp 1669390400
transform -1 0 26768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_93
timestamp 1669390400
transform -1 0 27440 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_94
timestamp 1669390400
transform -1 0 28112 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_95
timestamp 1669390400
transform -1 0 28784 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_96
timestamp 1669390400
transform -1 0 29456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_97
timestamp 1669390400
transform -1 0 30128 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_98
timestamp 1669390400
transform -1 0 3472 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_99
timestamp 1669390400
transform -1 0 5488 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_100
timestamp 1669390400
transform -1 0 7504 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_101
timestamp 1669390400
transform -1 0 9520 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_102
timestamp 1669390400
transform -1 0 11536 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_103
timestamp 1669390400
transform -1 0 13552 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_104
timestamp 1669390400
transform -1 0 15568 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_105
timestamp 1669390400
transform -1 0 17584 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_106
timestamp 1669390400
transform -1 0 19600 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_107
timestamp 1669390400
transform -1 0 22064 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_108
timestamp 1669390400
transform -1 0 23632 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_109
timestamp 1669390400
transform -1 0 25648 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_110
timestamp 1669390400
transform -1 0 27664 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_111
timestamp 1669390400
transform 1 0 28448 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_112
timestamp 1669390400
transform -1 0 31696 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_113
timestamp 1669390400
transform 1 0 32480 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_114
timestamp 1669390400
transform 1 0 34496 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_115
timestamp 1669390400
transform 1 0 36736 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_116
timestamp 1669390400
transform 1 0 36176 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_117
timestamp 1669390400
transform 1 0 40656 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_118
timestamp 1669390400
transform -1 0 46928 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_119
timestamp 1669390400
transform -1 0 46032 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_120
timestamp 1669390400
transform -1 0 48832 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_121
timestamp 1669390400
transform 1 0 48832 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_122
timestamp 1669390400
transform -1 0 52640 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_123
timestamp 1669390400
transform -1 0 60816 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_124
timestamp 1669390400
transform -1 0 60144 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_125
timestamp 1669390400
transform -1 0 60816 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_126
timestamp 1669390400
transform -1 0 60704 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_127
timestamp 1669390400
transform -1 0 63392 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_128
timestamp 1669390400
transform -1 0 64064 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_129
timestamp 1669390400
transform -1 0 65968 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_130
timestamp 1669390400
transform -1 0 67984 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_131
timestamp 1669390400
transform -1 0 70336 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_132
timestamp 1669390400
transform -1 0 72016 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_133
timestamp 1669390400
transform -1 0 74256 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_134
timestamp 1669390400
transform -1 0 76048 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_135
timestamp 1669390400
transform -1 0 78288 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_136
timestamp 1669390400
transform -1 0 6160 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_137
timestamp 1669390400
transform -1 0 8176 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_138
timestamp 1669390400
transform -1 0 10192 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_139
timestamp 1669390400
transform 1 0 34160 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_140
timestamp 1669390400
transform 1 0 37296 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_141
timestamp 1669390400
transform -1 0 47600 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_142
timestamp 1669390400
transform -1 0 47376 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_143
timestamp 1669390400
transform -1 0 48496 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_144
timestamp 1669390400
transform -1 0 50512 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_145
timestamp 1669390400
transform -1 0 60144 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_146
timestamp 1669390400
transform -1 0 60816 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_147
timestamp 1669390400
transform -1 0 62048 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_148
timestamp 1669390400
transform -1 0 62720 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_149
timestamp 1669390400
transform -1 0 62496 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_150
timestamp 1669390400
transform -1 0 63168 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_151
timestamp 1669390400
transform -1 0 64736 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_152
timestamp 1669390400
transform -1 0 66640 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_153
timestamp 1669390400
transform -1 0 70224 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_154
timestamp 1669390400
transform -1 0 71008 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_155
timestamp 1669390400
transform -1 0 72688 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_156
timestamp 1669390400
transform -1 0 74704 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_157
timestamp 1669390400
transform -1 0 76720 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_158
timestamp 1669390400
transform 1 0 77840 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_159
timestamp 1669390400
transform -1 0 73584 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_160
timestamp 1669390400
transform -1 0 74704 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_161
timestamp 1669390400
transform -1 0 74256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_162
timestamp 1669390400
transform -1 0 30800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_163
timestamp 1669390400
transform -1 0 31472 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_164
timestamp 1669390400
transform -1 0 32144 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_165
timestamp 1669390400
transform -1 0 32816 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_166
timestamp 1669390400
transform -1 0 33488 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_167
timestamp 1669390400
transform -1 0 34160 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_168
timestamp 1669390400
transform -1 0 34832 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_169
timestamp 1669390400
transform -1 0 35504 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_170
timestamp 1669390400
transform -1 0 36176 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_171
timestamp 1669390400
transform -1 0 36848 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_172
timestamp 1669390400
transform -1 0 37520 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_173
timestamp 1669390400
transform -1 0 38192 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_174
timestamp 1669390400
transform -1 0 38864 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_175
timestamp 1669390400
transform -1 0 39536 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_176
timestamp 1669390400
transform -1 0 40208 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_177
timestamp 1669390400
transform -1 0 40880 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_178
timestamp 1669390400
transform -1 0 42000 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_179
timestamp 1669390400
transform -1 0 42672 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_180
timestamp 1669390400
transform -1 0 43344 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_181
timestamp 1669390400
transform -1 0 44016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_182
timestamp 1669390400
transform -1 0 44688 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_183
timestamp 1669390400
transform -1 0 45360 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_184
timestamp 1669390400
transform -1 0 46032 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_185
timestamp 1669390400
transform -1 0 46704 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_186
timestamp 1669390400
transform -1 0 47376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_187
timestamp 1669390400
transform -1 0 48048 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_188
timestamp 1669390400
transform -1 0 48720 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_189
timestamp 1669390400
transform -1 0 49392 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_190
timestamp 1669390400
transform -1 0 50064 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_191
timestamp 1669390400
transform -1 0 50736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_192
timestamp 1669390400
transform -1 0 51408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_193
timestamp 1669390400
transform -1 0 52080 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_194
timestamp 1669390400
transform -1 0 52752 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_195
timestamp 1669390400
transform -1 0 53424 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_196
timestamp 1669390400
transform -1 0 54096 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  macro_tap_197
timestamp 1669390400
transform -1 0 54768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output22 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 5264 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output23
timestamp 1669390400
transform -1 0 25424 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output24
timestamp 1669390400
transform -1 0 27440 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output25
timestamp 1669390400
transform 1 0 27888 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output26
timestamp 1669390400
transform 1 0 29904 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output27
timestamp 1669390400
transform 1 0 31920 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output28
timestamp 1669390400
transform 1 0 33936 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output29
timestamp 1669390400
transform 1 0 35952 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output30
timestamp 1669390400
transform 1 0 37968 0 1 75264
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output31
timestamp 1669390400
transform -1 0 13328 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output32
timestamp 1669390400
transform -1 0 15344 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output33
timestamp 1669390400
transform -1 0 17360 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output34
timestamp 1669390400
transform -1 0 19376 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output35
timestamp 1669390400
transform -1 0 21168 0 -1 76832
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output36
timestamp 1669390400
transform -1 0 23408 0 -1 76832
box -86 -86 1654 870
<< labels >>
flabel metal2 s 1568 79200 1680 80000 0 FreeSans 448 90 0 0 io_active
port 0 nsew signal input
flabel metal2 s 2240 79200 2352 80000 0 FreeSans 448 90 0 0 io_in[0]
port 1 nsew signal input
flabel metal2 s 22400 79200 22512 80000 0 FreeSans 448 90 0 0 io_in[10]
port 2 nsew signal input
flabel metal2 s 24416 79200 24528 80000 0 FreeSans 448 90 0 0 io_in[11]
port 3 nsew signal input
flabel metal2 s 26432 79200 26544 80000 0 FreeSans 448 90 0 0 io_in[12]
port 4 nsew signal input
flabel metal2 s 28448 79200 28560 80000 0 FreeSans 448 90 0 0 io_in[13]
port 5 nsew signal input
flabel metal2 s 30464 79200 30576 80000 0 FreeSans 448 90 0 0 io_in[14]
port 6 nsew signal input
flabel metal2 s 32480 79200 32592 80000 0 FreeSans 448 90 0 0 io_in[15]
port 7 nsew signal input
flabel metal2 s 34496 79200 34608 80000 0 FreeSans 448 90 0 0 io_in[16]
port 8 nsew signal input
flabel metal2 s 36512 79200 36624 80000 0 FreeSans 448 90 0 0 io_in[17]
port 9 nsew signal input
flabel metal2 s 38528 79200 38640 80000 0 FreeSans 448 90 0 0 io_in[18]
port 10 nsew signal input
flabel metal2 s 40544 79200 40656 80000 0 FreeSans 448 90 0 0 io_in[19]
port 11 nsew signal input
flabel metal2 s 4256 79200 4368 80000 0 FreeSans 448 90 0 0 io_in[1]
port 12 nsew signal input
flabel metal2 s 42560 79200 42672 80000 0 FreeSans 448 90 0 0 io_in[20]
port 13 nsew signal input
flabel metal2 s 44576 79200 44688 80000 0 FreeSans 448 90 0 0 io_in[21]
port 14 nsew signal input
flabel metal2 s 46592 79200 46704 80000 0 FreeSans 448 90 0 0 io_in[22]
port 15 nsew signal input
flabel metal2 s 48608 79200 48720 80000 0 FreeSans 448 90 0 0 io_in[23]
port 16 nsew signal input
flabel metal2 s 50624 79200 50736 80000 0 FreeSans 448 90 0 0 io_in[24]
port 17 nsew signal input
flabel metal2 s 52640 79200 52752 80000 0 FreeSans 448 90 0 0 io_in[25]
port 18 nsew signal input
flabel metal2 s 54656 79200 54768 80000 0 FreeSans 448 90 0 0 io_in[26]
port 19 nsew signal input
flabel metal2 s 56672 79200 56784 80000 0 FreeSans 448 90 0 0 io_in[27]
port 20 nsew signal input
flabel metal2 s 58688 79200 58800 80000 0 FreeSans 448 90 0 0 io_in[28]
port 21 nsew signal input
flabel metal2 s 60704 79200 60816 80000 0 FreeSans 448 90 0 0 io_in[29]
port 22 nsew signal input
flabel metal2 s 6272 79200 6384 80000 0 FreeSans 448 90 0 0 io_in[2]
port 23 nsew signal input
flabel metal2 s 62720 79200 62832 80000 0 FreeSans 448 90 0 0 io_in[30]
port 24 nsew signal input
flabel metal2 s 64736 79200 64848 80000 0 FreeSans 448 90 0 0 io_in[31]
port 25 nsew signal input
flabel metal2 s 66752 79200 66864 80000 0 FreeSans 448 90 0 0 io_in[32]
port 26 nsew signal input
flabel metal2 s 68768 79200 68880 80000 0 FreeSans 448 90 0 0 io_in[33]
port 27 nsew signal input
flabel metal2 s 70784 79200 70896 80000 0 FreeSans 448 90 0 0 io_in[34]
port 28 nsew signal input
flabel metal2 s 72800 79200 72912 80000 0 FreeSans 448 90 0 0 io_in[35]
port 29 nsew signal input
flabel metal2 s 74816 79200 74928 80000 0 FreeSans 448 90 0 0 io_in[36]
port 30 nsew signal input
flabel metal2 s 76832 79200 76944 80000 0 FreeSans 448 90 0 0 io_in[37]
port 31 nsew signal input
flabel metal2 s 8288 79200 8400 80000 0 FreeSans 448 90 0 0 io_in[3]
port 32 nsew signal input
flabel metal2 s 10304 79200 10416 80000 0 FreeSans 448 90 0 0 io_in[4]
port 33 nsew signal input
flabel metal2 s 12320 79200 12432 80000 0 FreeSans 448 90 0 0 io_in[5]
port 34 nsew signal input
flabel metal2 s 14336 79200 14448 80000 0 FreeSans 448 90 0 0 io_in[6]
port 35 nsew signal input
flabel metal2 s 16352 79200 16464 80000 0 FreeSans 448 90 0 0 io_in[7]
port 36 nsew signal input
flabel metal2 s 18368 79200 18480 80000 0 FreeSans 448 90 0 0 io_in[8]
port 37 nsew signal input
flabel metal2 s 20384 79200 20496 80000 0 FreeSans 448 90 0 0 io_in[9]
port 38 nsew signal input
flabel metal2 s 2912 79200 3024 80000 0 FreeSans 448 90 0 0 io_oeb[0]
port 39 nsew signal tristate
flabel metal2 s 23072 79200 23184 80000 0 FreeSans 448 90 0 0 io_oeb[10]
port 40 nsew signal tristate
flabel metal2 s 25088 79200 25200 80000 0 FreeSans 448 90 0 0 io_oeb[11]
port 41 nsew signal tristate
flabel metal2 s 27104 79200 27216 80000 0 FreeSans 448 90 0 0 io_oeb[12]
port 42 nsew signal tristate
flabel metal2 s 29120 79200 29232 80000 0 FreeSans 448 90 0 0 io_oeb[13]
port 43 nsew signal tristate
flabel metal2 s 31136 79200 31248 80000 0 FreeSans 448 90 0 0 io_oeb[14]
port 44 nsew signal tristate
flabel metal2 s 33152 79200 33264 80000 0 FreeSans 448 90 0 0 io_oeb[15]
port 45 nsew signal tristate
flabel metal2 s 35168 79200 35280 80000 0 FreeSans 448 90 0 0 io_oeb[16]
port 46 nsew signal tristate
flabel metal2 s 37184 79200 37296 80000 0 FreeSans 448 90 0 0 io_oeb[17]
port 47 nsew signal tristate
flabel metal2 s 39200 79200 39312 80000 0 FreeSans 448 90 0 0 io_oeb[18]
port 48 nsew signal tristate
flabel metal2 s 41216 79200 41328 80000 0 FreeSans 448 90 0 0 io_oeb[19]
port 49 nsew signal tristate
flabel metal2 s 4928 79200 5040 80000 0 FreeSans 448 90 0 0 io_oeb[1]
port 50 nsew signal tristate
flabel metal2 s 43232 79200 43344 80000 0 FreeSans 448 90 0 0 io_oeb[20]
port 51 nsew signal tristate
flabel metal2 s 45248 79200 45360 80000 0 FreeSans 448 90 0 0 io_oeb[21]
port 52 nsew signal tristate
flabel metal2 s 47264 79200 47376 80000 0 FreeSans 448 90 0 0 io_oeb[22]
port 53 nsew signal tristate
flabel metal2 s 49280 79200 49392 80000 0 FreeSans 448 90 0 0 io_oeb[23]
port 54 nsew signal tristate
flabel metal2 s 51296 79200 51408 80000 0 FreeSans 448 90 0 0 io_oeb[24]
port 55 nsew signal tristate
flabel metal2 s 53312 79200 53424 80000 0 FreeSans 448 90 0 0 io_oeb[25]
port 56 nsew signal tristate
flabel metal2 s 55328 79200 55440 80000 0 FreeSans 448 90 0 0 io_oeb[26]
port 57 nsew signal tristate
flabel metal2 s 57344 79200 57456 80000 0 FreeSans 448 90 0 0 io_oeb[27]
port 58 nsew signal tristate
flabel metal2 s 59360 79200 59472 80000 0 FreeSans 448 90 0 0 io_oeb[28]
port 59 nsew signal tristate
flabel metal2 s 61376 79200 61488 80000 0 FreeSans 448 90 0 0 io_oeb[29]
port 60 nsew signal tristate
flabel metal2 s 6944 79200 7056 80000 0 FreeSans 448 90 0 0 io_oeb[2]
port 61 nsew signal tristate
flabel metal2 s 63392 79200 63504 80000 0 FreeSans 448 90 0 0 io_oeb[30]
port 62 nsew signal tristate
flabel metal2 s 65408 79200 65520 80000 0 FreeSans 448 90 0 0 io_oeb[31]
port 63 nsew signal tristate
flabel metal2 s 67424 79200 67536 80000 0 FreeSans 448 90 0 0 io_oeb[32]
port 64 nsew signal tristate
flabel metal2 s 69440 79200 69552 80000 0 FreeSans 448 90 0 0 io_oeb[33]
port 65 nsew signal tristate
flabel metal2 s 71456 79200 71568 80000 0 FreeSans 448 90 0 0 io_oeb[34]
port 66 nsew signal tristate
flabel metal2 s 73472 79200 73584 80000 0 FreeSans 448 90 0 0 io_oeb[35]
port 67 nsew signal tristate
flabel metal2 s 75488 79200 75600 80000 0 FreeSans 448 90 0 0 io_oeb[36]
port 68 nsew signal tristate
flabel metal2 s 77504 79200 77616 80000 0 FreeSans 448 90 0 0 io_oeb[37]
port 69 nsew signal tristate
flabel metal2 s 8960 79200 9072 80000 0 FreeSans 448 90 0 0 io_oeb[3]
port 70 nsew signal tristate
flabel metal2 s 10976 79200 11088 80000 0 FreeSans 448 90 0 0 io_oeb[4]
port 71 nsew signal tristate
flabel metal2 s 12992 79200 13104 80000 0 FreeSans 448 90 0 0 io_oeb[5]
port 72 nsew signal tristate
flabel metal2 s 15008 79200 15120 80000 0 FreeSans 448 90 0 0 io_oeb[6]
port 73 nsew signal tristate
flabel metal2 s 17024 79200 17136 80000 0 FreeSans 448 90 0 0 io_oeb[7]
port 74 nsew signal tristate
flabel metal2 s 19040 79200 19152 80000 0 FreeSans 448 90 0 0 io_oeb[8]
port 75 nsew signal tristate
flabel metal2 s 21056 79200 21168 80000 0 FreeSans 448 90 0 0 io_oeb[9]
port 76 nsew signal tristate
flabel metal2 s 3584 79200 3696 80000 0 FreeSans 448 90 0 0 io_out[0]
port 77 nsew signal tristate
flabel metal2 s 23744 79200 23856 80000 0 FreeSans 448 90 0 0 io_out[10]
port 78 nsew signal tristate
flabel metal2 s 25760 79200 25872 80000 0 FreeSans 448 90 0 0 io_out[11]
port 79 nsew signal tristate
flabel metal2 s 27776 79200 27888 80000 0 FreeSans 448 90 0 0 io_out[12]
port 80 nsew signal tristate
flabel metal2 s 29792 79200 29904 80000 0 FreeSans 448 90 0 0 io_out[13]
port 81 nsew signal tristate
flabel metal2 s 31808 79200 31920 80000 0 FreeSans 448 90 0 0 io_out[14]
port 82 nsew signal tristate
flabel metal2 s 33824 79200 33936 80000 0 FreeSans 448 90 0 0 io_out[15]
port 83 nsew signal tristate
flabel metal2 s 35840 79200 35952 80000 0 FreeSans 448 90 0 0 io_out[16]
port 84 nsew signal tristate
flabel metal2 s 37856 79200 37968 80000 0 FreeSans 448 90 0 0 io_out[17]
port 85 nsew signal tristate
flabel metal2 s 39872 79200 39984 80000 0 FreeSans 448 90 0 0 io_out[18]
port 86 nsew signal tristate
flabel metal2 s 41888 79200 42000 80000 0 FreeSans 448 90 0 0 io_out[19]
port 87 nsew signal tristate
flabel metal2 s 5600 79200 5712 80000 0 FreeSans 448 90 0 0 io_out[1]
port 88 nsew signal tristate
flabel metal2 s 43904 79200 44016 80000 0 FreeSans 448 90 0 0 io_out[20]
port 89 nsew signal tristate
flabel metal2 s 45920 79200 46032 80000 0 FreeSans 448 90 0 0 io_out[21]
port 90 nsew signal tristate
flabel metal2 s 47936 79200 48048 80000 0 FreeSans 448 90 0 0 io_out[22]
port 91 nsew signal tristate
flabel metal2 s 49952 79200 50064 80000 0 FreeSans 448 90 0 0 io_out[23]
port 92 nsew signal tristate
flabel metal2 s 51968 79200 52080 80000 0 FreeSans 448 90 0 0 io_out[24]
port 93 nsew signal tristate
flabel metal2 s 53984 79200 54096 80000 0 FreeSans 448 90 0 0 io_out[25]
port 94 nsew signal tristate
flabel metal2 s 56000 79200 56112 80000 0 FreeSans 448 90 0 0 io_out[26]
port 95 nsew signal tristate
flabel metal2 s 58016 79200 58128 80000 0 FreeSans 448 90 0 0 io_out[27]
port 96 nsew signal tristate
flabel metal2 s 60032 79200 60144 80000 0 FreeSans 448 90 0 0 io_out[28]
port 97 nsew signal tristate
flabel metal2 s 62048 79200 62160 80000 0 FreeSans 448 90 0 0 io_out[29]
port 98 nsew signal tristate
flabel metal2 s 7616 79200 7728 80000 0 FreeSans 448 90 0 0 io_out[2]
port 99 nsew signal tristate
flabel metal2 s 64064 79200 64176 80000 0 FreeSans 448 90 0 0 io_out[30]
port 100 nsew signal tristate
flabel metal2 s 66080 79200 66192 80000 0 FreeSans 448 90 0 0 io_out[31]
port 101 nsew signal tristate
flabel metal2 s 68096 79200 68208 80000 0 FreeSans 448 90 0 0 io_out[32]
port 102 nsew signal tristate
flabel metal2 s 70112 79200 70224 80000 0 FreeSans 448 90 0 0 io_out[33]
port 103 nsew signal tristate
flabel metal2 s 72128 79200 72240 80000 0 FreeSans 448 90 0 0 io_out[34]
port 104 nsew signal tristate
flabel metal2 s 74144 79200 74256 80000 0 FreeSans 448 90 0 0 io_out[35]
port 105 nsew signal tristate
flabel metal2 s 76160 79200 76272 80000 0 FreeSans 448 90 0 0 io_out[36]
port 106 nsew signal tristate
flabel metal2 s 78176 79200 78288 80000 0 FreeSans 448 90 0 0 io_out[37]
port 107 nsew signal tristate
flabel metal2 s 9632 79200 9744 80000 0 FreeSans 448 90 0 0 io_out[3]
port 108 nsew signal tristate
flabel metal2 s 11648 79200 11760 80000 0 FreeSans 448 90 0 0 io_out[4]
port 109 nsew signal tristate
flabel metal2 s 13664 79200 13776 80000 0 FreeSans 448 90 0 0 io_out[5]
port 110 nsew signal tristate
flabel metal2 s 15680 79200 15792 80000 0 FreeSans 448 90 0 0 io_out[6]
port 111 nsew signal tristate
flabel metal2 s 17696 79200 17808 80000 0 FreeSans 448 90 0 0 io_out[7]
port 112 nsew signal tristate
flabel metal2 s 19712 79200 19824 80000 0 FreeSans 448 90 0 0 io_out[8]
port 113 nsew signal tristate
flabel metal2 s 21728 79200 21840 80000 0 FreeSans 448 90 0 0 io_out[9]
port 114 nsew signal tristate
flabel metal2 s 73024 0 73136 800 0 FreeSans 448 90 0 0 irq[0]
port 115 nsew signal tristate
flabel metal2 s 73248 0 73360 800 0 FreeSans 448 90 0 0 irq[1]
port 116 nsew signal tristate
flabel metal2 s 73472 0 73584 800 0 FreeSans 448 90 0 0 irq[2]
port 117 nsew signal tristate
flabel metal2 s 30016 0 30128 800 0 FreeSans 448 90 0 0 la_data_in[0]
port 118 nsew signal input
flabel metal2 s 36736 0 36848 800 0 FreeSans 448 90 0 0 la_data_in[10]
port 119 nsew signal input
flabel metal2 s 37408 0 37520 800 0 FreeSans 448 90 0 0 la_data_in[11]
port 120 nsew signal input
flabel metal2 s 38080 0 38192 800 0 FreeSans 448 90 0 0 la_data_in[12]
port 121 nsew signal input
flabel metal2 s 38752 0 38864 800 0 FreeSans 448 90 0 0 la_data_in[13]
port 122 nsew signal input
flabel metal2 s 39424 0 39536 800 0 FreeSans 448 90 0 0 la_data_in[14]
port 123 nsew signal input
flabel metal2 s 40096 0 40208 800 0 FreeSans 448 90 0 0 la_data_in[15]
port 124 nsew signal input
flabel metal2 s 40768 0 40880 800 0 FreeSans 448 90 0 0 la_data_in[16]
port 125 nsew signal input
flabel metal2 s 41440 0 41552 800 0 FreeSans 448 90 0 0 la_data_in[17]
port 126 nsew signal input
flabel metal2 s 42112 0 42224 800 0 FreeSans 448 90 0 0 la_data_in[18]
port 127 nsew signal input
flabel metal2 s 42784 0 42896 800 0 FreeSans 448 90 0 0 la_data_in[19]
port 128 nsew signal input
flabel metal2 s 30688 0 30800 800 0 FreeSans 448 90 0 0 la_data_in[1]
port 129 nsew signal input
flabel metal2 s 43456 0 43568 800 0 FreeSans 448 90 0 0 la_data_in[20]
port 130 nsew signal input
flabel metal2 s 44128 0 44240 800 0 FreeSans 448 90 0 0 la_data_in[21]
port 131 nsew signal input
flabel metal2 s 44800 0 44912 800 0 FreeSans 448 90 0 0 la_data_in[22]
port 132 nsew signal input
flabel metal2 s 45472 0 45584 800 0 FreeSans 448 90 0 0 la_data_in[23]
port 133 nsew signal input
flabel metal2 s 46144 0 46256 800 0 FreeSans 448 90 0 0 la_data_in[24]
port 134 nsew signal input
flabel metal2 s 46816 0 46928 800 0 FreeSans 448 90 0 0 la_data_in[25]
port 135 nsew signal input
flabel metal2 s 47488 0 47600 800 0 FreeSans 448 90 0 0 la_data_in[26]
port 136 nsew signal input
flabel metal2 s 48160 0 48272 800 0 FreeSans 448 90 0 0 la_data_in[27]
port 137 nsew signal input
flabel metal2 s 48832 0 48944 800 0 FreeSans 448 90 0 0 la_data_in[28]
port 138 nsew signal input
flabel metal2 s 49504 0 49616 800 0 FreeSans 448 90 0 0 la_data_in[29]
port 139 nsew signal input
flabel metal2 s 31360 0 31472 800 0 FreeSans 448 90 0 0 la_data_in[2]
port 140 nsew signal input
flabel metal2 s 50176 0 50288 800 0 FreeSans 448 90 0 0 la_data_in[30]
port 141 nsew signal input
flabel metal2 s 50848 0 50960 800 0 FreeSans 448 90 0 0 la_data_in[31]
port 142 nsew signal input
flabel metal2 s 51520 0 51632 800 0 FreeSans 448 90 0 0 la_data_in[32]
port 143 nsew signal input
flabel metal2 s 52192 0 52304 800 0 FreeSans 448 90 0 0 la_data_in[33]
port 144 nsew signal input
flabel metal2 s 52864 0 52976 800 0 FreeSans 448 90 0 0 la_data_in[34]
port 145 nsew signal input
flabel metal2 s 53536 0 53648 800 0 FreeSans 448 90 0 0 la_data_in[35]
port 146 nsew signal input
flabel metal2 s 54208 0 54320 800 0 FreeSans 448 90 0 0 la_data_in[36]
port 147 nsew signal input
flabel metal2 s 54880 0 54992 800 0 FreeSans 448 90 0 0 la_data_in[37]
port 148 nsew signal input
flabel metal2 s 55552 0 55664 800 0 FreeSans 448 90 0 0 la_data_in[38]
port 149 nsew signal input
flabel metal2 s 56224 0 56336 800 0 FreeSans 448 90 0 0 la_data_in[39]
port 150 nsew signal input
flabel metal2 s 32032 0 32144 800 0 FreeSans 448 90 0 0 la_data_in[3]
port 151 nsew signal input
flabel metal2 s 56896 0 57008 800 0 FreeSans 448 90 0 0 la_data_in[40]
port 152 nsew signal input
flabel metal2 s 57568 0 57680 800 0 FreeSans 448 90 0 0 la_data_in[41]
port 153 nsew signal input
flabel metal2 s 58240 0 58352 800 0 FreeSans 448 90 0 0 la_data_in[42]
port 154 nsew signal input
flabel metal2 s 58912 0 59024 800 0 FreeSans 448 90 0 0 la_data_in[43]
port 155 nsew signal input
flabel metal2 s 59584 0 59696 800 0 FreeSans 448 90 0 0 la_data_in[44]
port 156 nsew signal input
flabel metal2 s 60256 0 60368 800 0 FreeSans 448 90 0 0 la_data_in[45]
port 157 nsew signal input
flabel metal2 s 60928 0 61040 800 0 FreeSans 448 90 0 0 la_data_in[46]
port 158 nsew signal input
flabel metal2 s 61600 0 61712 800 0 FreeSans 448 90 0 0 la_data_in[47]
port 159 nsew signal input
flabel metal2 s 62272 0 62384 800 0 FreeSans 448 90 0 0 la_data_in[48]
port 160 nsew signal input
flabel metal2 s 62944 0 63056 800 0 FreeSans 448 90 0 0 la_data_in[49]
port 161 nsew signal input
flabel metal2 s 32704 0 32816 800 0 FreeSans 448 90 0 0 la_data_in[4]
port 162 nsew signal input
flabel metal2 s 63616 0 63728 800 0 FreeSans 448 90 0 0 la_data_in[50]
port 163 nsew signal input
flabel metal2 s 64288 0 64400 800 0 FreeSans 448 90 0 0 la_data_in[51]
port 164 nsew signal input
flabel metal2 s 64960 0 65072 800 0 FreeSans 448 90 0 0 la_data_in[52]
port 165 nsew signal input
flabel metal2 s 65632 0 65744 800 0 FreeSans 448 90 0 0 la_data_in[53]
port 166 nsew signal input
flabel metal2 s 66304 0 66416 800 0 FreeSans 448 90 0 0 la_data_in[54]
port 167 nsew signal input
flabel metal2 s 66976 0 67088 800 0 FreeSans 448 90 0 0 la_data_in[55]
port 168 nsew signal input
flabel metal2 s 67648 0 67760 800 0 FreeSans 448 90 0 0 la_data_in[56]
port 169 nsew signal input
flabel metal2 s 68320 0 68432 800 0 FreeSans 448 90 0 0 la_data_in[57]
port 170 nsew signal input
flabel metal2 s 68992 0 69104 800 0 FreeSans 448 90 0 0 la_data_in[58]
port 171 nsew signal input
flabel metal2 s 69664 0 69776 800 0 FreeSans 448 90 0 0 la_data_in[59]
port 172 nsew signal input
flabel metal2 s 33376 0 33488 800 0 FreeSans 448 90 0 0 la_data_in[5]
port 173 nsew signal input
flabel metal2 s 70336 0 70448 800 0 FreeSans 448 90 0 0 la_data_in[60]
port 174 nsew signal input
flabel metal2 s 71008 0 71120 800 0 FreeSans 448 90 0 0 la_data_in[61]
port 175 nsew signal input
flabel metal2 s 71680 0 71792 800 0 FreeSans 448 90 0 0 la_data_in[62]
port 176 nsew signal input
flabel metal2 s 72352 0 72464 800 0 FreeSans 448 90 0 0 la_data_in[63]
port 177 nsew signal input
flabel metal2 s 34048 0 34160 800 0 FreeSans 448 90 0 0 la_data_in[6]
port 178 nsew signal input
flabel metal2 s 34720 0 34832 800 0 FreeSans 448 90 0 0 la_data_in[7]
port 179 nsew signal input
flabel metal2 s 35392 0 35504 800 0 FreeSans 448 90 0 0 la_data_in[8]
port 180 nsew signal input
flabel metal2 s 36064 0 36176 800 0 FreeSans 448 90 0 0 la_data_in[9]
port 181 nsew signal input
flabel metal2 s 30240 0 30352 800 0 FreeSans 448 90 0 0 la_data_out[0]
port 182 nsew signal tristate
flabel metal2 s 36960 0 37072 800 0 FreeSans 448 90 0 0 la_data_out[10]
port 183 nsew signal tristate
flabel metal2 s 37632 0 37744 800 0 FreeSans 448 90 0 0 la_data_out[11]
port 184 nsew signal tristate
flabel metal2 s 38304 0 38416 800 0 FreeSans 448 90 0 0 la_data_out[12]
port 185 nsew signal tristate
flabel metal2 s 38976 0 39088 800 0 FreeSans 448 90 0 0 la_data_out[13]
port 186 nsew signal tristate
flabel metal2 s 39648 0 39760 800 0 FreeSans 448 90 0 0 la_data_out[14]
port 187 nsew signal tristate
flabel metal2 s 40320 0 40432 800 0 FreeSans 448 90 0 0 la_data_out[15]
port 188 nsew signal tristate
flabel metal2 s 40992 0 41104 800 0 FreeSans 448 90 0 0 la_data_out[16]
port 189 nsew signal tristate
flabel metal2 s 41664 0 41776 800 0 FreeSans 448 90 0 0 la_data_out[17]
port 190 nsew signal tristate
flabel metal2 s 42336 0 42448 800 0 FreeSans 448 90 0 0 la_data_out[18]
port 191 nsew signal tristate
flabel metal2 s 43008 0 43120 800 0 FreeSans 448 90 0 0 la_data_out[19]
port 192 nsew signal tristate
flabel metal2 s 30912 0 31024 800 0 FreeSans 448 90 0 0 la_data_out[1]
port 193 nsew signal tristate
flabel metal2 s 43680 0 43792 800 0 FreeSans 448 90 0 0 la_data_out[20]
port 194 nsew signal tristate
flabel metal2 s 44352 0 44464 800 0 FreeSans 448 90 0 0 la_data_out[21]
port 195 nsew signal tristate
flabel metal2 s 45024 0 45136 800 0 FreeSans 448 90 0 0 la_data_out[22]
port 196 nsew signal tristate
flabel metal2 s 45696 0 45808 800 0 FreeSans 448 90 0 0 la_data_out[23]
port 197 nsew signal tristate
flabel metal2 s 46368 0 46480 800 0 FreeSans 448 90 0 0 la_data_out[24]
port 198 nsew signal tristate
flabel metal2 s 47040 0 47152 800 0 FreeSans 448 90 0 0 la_data_out[25]
port 199 nsew signal tristate
flabel metal2 s 47712 0 47824 800 0 FreeSans 448 90 0 0 la_data_out[26]
port 200 nsew signal tristate
flabel metal2 s 48384 0 48496 800 0 FreeSans 448 90 0 0 la_data_out[27]
port 201 nsew signal tristate
flabel metal2 s 49056 0 49168 800 0 FreeSans 448 90 0 0 la_data_out[28]
port 202 nsew signal tristate
flabel metal2 s 49728 0 49840 800 0 FreeSans 448 90 0 0 la_data_out[29]
port 203 nsew signal tristate
flabel metal2 s 31584 0 31696 800 0 FreeSans 448 90 0 0 la_data_out[2]
port 204 nsew signal tristate
flabel metal2 s 50400 0 50512 800 0 FreeSans 448 90 0 0 la_data_out[30]
port 205 nsew signal tristate
flabel metal2 s 51072 0 51184 800 0 FreeSans 448 90 0 0 la_data_out[31]
port 206 nsew signal tristate
flabel metal2 s 51744 0 51856 800 0 FreeSans 448 90 0 0 la_data_out[32]
port 207 nsew signal tristate
flabel metal2 s 52416 0 52528 800 0 FreeSans 448 90 0 0 la_data_out[33]
port 208 nsew signal tristate
flabel metal2 s 53088 0 53200 800 0 FreeSans 448 90 0 0 la_data_out[34]
port 209 nsew signal tristate
flabel metal2 s 53760 0 53872 800 0 FreeSans 448 90 0 0 la_data_out[35]
port 210 nsew signal tristate
flabel metal2 s 54432 0 54544 800 0 FreeSans 448 90 0 0 la_data_out[36]
port 211 nsew signal tristate
flabel metal2 s 55104 0 55216 800 0 FreeSans 448 90 0 0 la_data_out[37]
port 212 nsew signal tristate
flabel metal2 s 55776 0 55888 800 0 FreeSans 448 90 0 0 la_data_out[38]
port 213 nsew signal tristate
flabel metal2 s 56448 0 56560 800 0 FreeSans 448 90 0 0 la_data_out[39]
port 214 nsew signal tristate
flabel metal2 s 32256 0 32368 800 0 FreeSans 448 90 0 0 la_data_out[3]
port 215 nsew signal tristate
flabel metal2 s 57120 0 57232 800 0 FreeSans 448 90 0 0 la_data_out[40]
port 216 nsew signal tristate
flabel metal2 s 57792 0 57904 800 0 FreeSans 448 90 0 0 la_data_out[41]
port 217 nsew signal tristate
flabel metal2 s 58464 0 58576 800 0 FreeSans 448 90 0 0 la_data_out[42]
port 218 nsew signal tristate
flabel metal2 s 59136 0 59248 800 0 FreeSans 448 90 0 0 la_data_out[43]
port 219 nsew signal tristate
flabel metal2 s 59808 0 59920 800 0 FreeSans 448 90 0 0 la_data_out[44]
port 220 nsew signal tristate
flabel metal2 s 60480 0 60592 800 0 FreeSans 448 90 0 0 la_data_out[45]
port 221 nsew signal tristate
flabel metal2 s 61152 0 61264 800 0 FreeSans 448 90 0 0 la_data_out[46]
port 222 nsew signal tristate
flabel metal2 s 61824 0 61936 800 0 FreeSans 448 90 0 0 la_data_out[47]
port 223 nsew signal tristate
flabel metal2 s 62496 0 62608 800 0 FreeSans 448 90 0 0 la_data_out[48]
port 224 nsew signal tristate
flabel metal2 s 63168 0 63280 800 0 FreeSans 448 90 0 0 la_data_out[49]
port 225 nsew signal tristate
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 la_data_out[4]
port 226 nsew signal tristate
flabel metal2 s 63840 0 63952 800 0 FreeSans 448 90 0 0 la_data_out[50]
port 227 nsew signal tristate
flabel metal2 s 64512 0 64624 800 0 FreeSans 448 90 0 0 la_data_out[51]
port 228 nsew signal tristate
flabel metal2 s 65184 0 65296 800 0 FreeSans 448 90 0 0 la_data_out[52]
port 229 nsew signal tristate
flabel metal2 s 65856 0 65968 800 0 FreeSans 448 90 0 0 la_data_out[53]
port 230 nsew signal tristate
flabel metal2 s 66528 0 66640 800 0 FreeSans 448 90 0 0 la_data_out[54]
port 231 nsew signal tristate
flabel metal2 s 67200 0 67312 800 0 FreeSans 448 90 0 0 la_data_out[55]
port 232 nsew signal tristate
flabel metal2 s 67872 0 67984 800 0 FreeSans 448 90 0 0 la_data_out[56]
port 233 nsew signal tristate
flabel metal2 s 68544 0 68656 800 0 FreeSans 448 90 0 0 la_data_out[57]
port 234 nsew signal tristate
flabel metal2 s 69216 0 69328 800 0 FreeSans 448 90 0 0 la_data_out[58]
port 235 nsew signal tristate
flabel metal2 s 69888 0 70000 800 0 FreeSans 448 90 0 0 la_data_out[59]
port 236 nsew signal tristate
flabel metal2 s 33600 0 33712 800 0 FreeSans 448 90 0 0 la_data_out[5]
port 237 nsew signal tristate
flabel metal2 s 70560 0 70672 800 0 FreeSans 448 90 0 0 la_data_out[60]
port 238 nsew signal tristate
flabel metal2 s 71232 0 71344 800 0 FreeSans 448 90 0 0 la_data_out[61]
port 239 nsew signal tristate
flabel metal2 s 71904 0 72016 800 0 FreeSans 448 90 0 0 la_data_out[62]
port 240 nsew signal tristate
flabel metal2 s 72576 0 72688 800 0 FreeSans 448 90 0 0 la_data_out[63]
port 241 nsew signal tristate
flabel metal2 s 34272 0 34384 800 0 FreeSans 448 90 0 0 la_data_out[6]
port 242 nsew signal tristate
flabel metal2 s 34944 0 35056 800 0 FreeSans 448 90 0 0 la_data_out[7]
port 243 nsew signal tristate
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 la_data_out[8]
port 244 nsew signal tristate
flabel metal2 s 36288 0 36400 800 0 FreeSans 448 90 0 0 la_data_out[9]
port 245 nsew signal tristate
flabel metal2 s 30464 0 30576 800 0 FreeSans 448 90 0 0 la_oenb[0]
port 246 nsew signal input
flabel metal2 s 37184 0 37296 800 0 FreeSans 448 90 0 0 la_oenb[10]
port 247 nsew signal input
flabel metal2 s 37856 0 37968 800 0 FreeSans 448 90 0 0 la_oenb[11]
port 248 nsew signal input
flabel metal2 s 38528 0 38640 800 0 FreeSans 448 90 0 0 la_oenb[12]
port 249 nsew signal input
flabel metal2 s 39200 0 39312 800 0 FreeSans 448 90 0 0 la_oenb[13]
port 250 nsew signal input
flabel metal2 s 39872 0 39984 800 0 FreeSans 448 90 0 0 la_oenb[14]
port 251 nsew signal input
flabel metal2 s 40544 0 40656 800 0 FreeSans 448 90 0 0 la_oenb[15]
port 252 nsew signal input
flabel metal2 s 41216 0 41328 800 0 FreeSans 448 90 0 0 la_oenb[16]
port 253 nsew signal input
flabel metal2 s 41888 0 42000 800 0 FreeSans 448 90 0 0 la_oenb[17]
port 254 nsew signal input
flabel metal2 s 42560 0 42672 800 0 FreeSans 448 90 0 0 la_oenb[18]
port 255 nsew signal input
flabel metal2 s 43232 0 43344 800 0 FreeSans 448 90 0 0 la_oenb[19]
port 256 nsew signal input
flabel metal2 s 31136 0 31248 800 0 FreeSans 448 90 0 0 la_oenb[1]
port 257 nsew signal input
flabel metal2 s 43904 0 44016 800 0 FreeSans 448 90 0 0 la_oenb[20]
port 258 nsew signal input
flabel metal2 s 44576 0 44688 800 0 FreeSans 448 90 0 0 la_oenb[21]
port 259 nsew signal input
flabel metal2 s 45248 0 45360 800 0 FreeSans 448 90 0 0 la_oenb[22]
port 260 nsew signal input
flabel metal2 s 45920 0 46032 800 0 FreeSans 448 90 0 0 la_oenb[23]
port 261 nsew signal input
flabel metal2 s 46592 0 46704 800 0 FreeSans 448 90 0 0 la_oenb[24]
port 262 nsew signal input
flabel metal2 s 47264 0 47376 800 0 FreeSans 448 90 0 0 la_oenb[25]
port 263 nsew signal input
flabel metal2 s 47936 0 48048 800 0 FreeSans 448 90 0 0 la_oenb[26]
port 264 nsew signal input
flabel metal2 s 48608 0 48720 800 0 FreeSans 448 90 0 0 la_oenb[27]
port 265 nsew signal input
flabel metal2 s 49280 0 49392 800 0 FreeSans 448 90 0 0 la_oenb[28]
port 266 nsew signal input
flabel metal2 s 49952 0 50064 800 0 FreeSans 448 90 0 0 la_oenb[29]
port 267 nsew signal input
flabel metal2 s 31808 0 31920 800 0 FreeSans 448 90 0 0 la_oenb[2]
port 268 nsew signal input
flabel metal2 s 50624 0 50736 800 0 FreeSans 448 90 0 0 la_oenb[30]
port 269 nsew signal input
flabel metal2 s 51296 0 51408 800 0 FreeSans 448 90 0 0 la_oenb[31]
port 270 nsew signal input
flabel metal2 s 51968 0 52080 800 0 FreeSans 448 90 0 0 la_oenb[32]
port 271 nsew signal input
flabel metal2 s 52640 0 52752 800 0 FreeSans 448 90 0 0 la_oenb[33]
port 272 nsew signal input
flabel metal2 s 53312 0 53424 800 0 FreeSans 448 90 0 0 la_oenb[34]
port 273 nsew signal input
flabel metal2 s 53984 0 54096 800 0 FreeSans 448 90 0 0 la_oenb[35]
port 274 nsew signal input
flabel metal2 s 54656 0 54768 800 0 FreeSans 448 90 0 0 la_oenb[36]
port 275 nsew signal input
flabel metal2 s 55328 0 55440 800 0 FreeSans 448 90 0 0 la_oenb[37]
port 276 nsew signal input
flabel metal2 s 56000 0 56112 800 0 FreeSans 448 90 0 0 la_oenb[38]
port 277 nsew signal input
flabel metal2 s 56672 0 56784 800 0 FreeSans 448 90 0 0 la_oenb[39]
port 278 nsew signal input
flabel metal2 s 32480 0 32592 800 0 FreeSans 448 90 0 0 la_oenb[3]
port 279 nsew signal input
flabel metal2 s 57344 0 57456 800 0 FreeSans 448 90 0 0 la_oenb[40]
port 280 nsew signal input
flabel metal2 s 58016 0 58128 800 0 FreeSans 448 90 0 0 la_oenb[41]
port 281 nsew signal input
flabel metal2 s 58688 0 58800 800 0 FreeSans 448 90 0 0 la_oenb[42]
port 282 nsew signal input
flabel metal2 s 59360 0 59472 800 0 FreeSans 448 90 0 0 la_oenb[43]
port 283 nsew signal input
flabel metal2 s 60032 0 60144 800 0 FreeSans 448 90 0 0 la_oenb[44]
port 284 nsew signal input
flabel metal2 s 60704 0 60816 800 0 FreeSans 448 90 0 0 la_oenb[45]
port 285 nsew signal input
flabel metal2 s 61376 0 61488 800 0 FreeSans 448 90 0 0 la_oenb[46]
port 286 nsew signal input
flabel metal2 s 62048 0 62160 800 0 FreeSans 448 90 0 0 la_oenb[47]
port 287 nsew signal input
flabel metal2 s 62720 0 62832 800 0 FreeSans 448 90 0 0 la_oenb[48]
port 288 nsew signal input
flabel metal2 s 63392 0 63504 800 0 FreeSans 448 90 0 0 la_oenb[49]
port 289 nsew signal input
flabel metal2 s 33152 0 33264 800 0 FreeSans 448 90 0 0 la_oenb[4]
port 290 nsew signal input
flabel metal2 s 64064 0 64176 800 0 FreeSans 448 90 0 0 la_oenb[50]
port 291 nsew signal input
flabel metal2 s 64736 0 64848 800 0 FreeSans 448 90 0 0 la_oenb[51]
port 292 nsew signal input
flabel metal2 s 65408 0 65520 800 0 FreeSans 448 90 0 0 la_oenb[52]
port 293 nsew signal input
flabel metal2 s 66080 0 66192 800 0 FreeSans 448 90 0 0 la_oenb[53]
port 294 nsew signal input
flabel metal2 s 66752 0 66864 800 0 FreeSans 448 90 0 0 la_oenb[54]
port 295 nsew signal input
flabel metal2 s 67424 0 67536 800 0 FreeSans 448 90 0 0 la_oenb[55]
port 296 nsew signal input
flabel metal2 s 68096 0 68208 800 0 FreeSans 448 90 0 0 la_oenb[56]
port 297 nsew signal input
flabel metal2 s 68768 0 68880 800 0 FreeSans 448 90 0 0 la_oenb[57]
port 298 nsew signal input
flabel metal2 s 69440 0 69552 800 0 FreeSans 448 90 0 0 la_oenb[58]
port 299 nsew signal input
flabel metal2 s 70112 0 70224 800 0 FreeSans 448 90 0 0 la_oenb[59]
port 300 nsew signal input
flabel metal2 s 33824 0 33936 800 0 FreeSans 448 90 0 0 la_oenb[5]
port 301 nsew signal input
flabel metal2 s 70784 0 70896 800 0 FreeSans 448 90 0 0 la_oenb[60]
port 302 nsew signal input
flabel metal2 s 71456 0 71568 800 0 FreeSans 448 90 0 0 la_oenb[61]
port 303 nsew signal input
flabel metal2 s 72128 0 72240 800 0 FreeSans 448 90 0 0 la_oenb[62]
port 304 nsew signal input
flabel metal2 s 72800 0 72912 800 0 FreeSans 448 90 0 0 la_oenb[63]
port 305 nsew signal input
flabel metal2 s 34496 0 34608 800 0 FreeSans 448 90 0 0 la_oenb[6]
port 306 nsew signal input
flabel metal2 s 35168 0 35280 800 0 FreeSans 448 90 0 0 la_oenb[7]
port 307 nsew signal input
flabel metal2 s 35840 0 35952 800 0 FreeSans 448 90 0 0 la_oenb[8]
port 308 nsew signal input
flabel metal2 s 36512 0 36624 800 0 FreeSans 448 90 0 0 la_oenb[9]
port 309 nsew signal input
flabel metal4 s 4448 3076 4768 76892 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 35168 3076 35488 76892 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 65888 3076 66208 76892 0 FreeSans 1280 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 19808 3076 20128 76892 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 76892 0 FreeSans 1280 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 6272 0 6384 800 0 FreeSans 448 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 6496 0 6608 800 0 FreeSans 448 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 7616 0 7728 800 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 15232 0 15344 800 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 15904 0 16016 800 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 16576 0 16688 800 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 17248 0 17360 800 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 17920 0 18032 800 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 18592 0 18704 800 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 19264 0 19376 800 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 19936 0 20048 800 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 20608 0 20720 800 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 21280 0 21392 800 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 8512 0 8624 800 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 21952 0 22064 800 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 22624 0 22736 800 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 23296 0 23408 800 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 23968 0 24080 800 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 24640 0 24752 800 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 25312 0 25424 800 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 25984 0 26096 800 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 26656 0 26768 800 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 27328 0 27440 800 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 28000 0 28112 800 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 28672 0 28784 800 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 29344 0 29456 800 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 10304 0 10416 800 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 11200 0 11312 800 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 11872 0 11984 800 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 12544 0 12656 800 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 13216 0 13328 800 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 13888 0 14000 800 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 14560 0 14672 800 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 6944 0 7056 800 0 FreeSans 448 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 7840 0 7952 800 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 21504 0 21616 800 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 27552 0 27664 800 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 28224 0 28336 800 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 9632 0 9744 800 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 10528 0 10640 800 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 11424 0 11536 800 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 12768 0 12880 800 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 14112 0 14224 800 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 15680 0 15792 800 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 16352 0 16464 800 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 17024 0 17136 800 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 17696 0 17808 800 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 18368 0 18480 800 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 19040 0 19152 800 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 19712 0 19824 800 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 20384 0 20496 800 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 21056 0 21168 800 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 21728 0 21840 800 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 8960 0 9072 800 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 22400 0 22512 800 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 23072 0 23184 800 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 23744 0 23856 800 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 24416 0 24528 800 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 25088 0 25200 800 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 25760 0 25872 800 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 26432 0 26544 800 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 27104 0 27216 800 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 27776 0 27888 800 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 28448 0 28560 800 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 9856 0 9968 800 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 29120 0 29232 800 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 29792 0 29904 800 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 11648 0 11760 800 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 12320 0 12432 800 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 12992 0 13104 800 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 13664 0 13776 800 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 14336 0 14448 800 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 15008 0 15120 800 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 8288 0 8400 800 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 9184 0 9296 800 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 10976 0 11088 800 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 7168 0 7280 800 0 FreeSans 448 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel metal1 39984 76048 39984 76048 0 vdd
rlabel metal1 39984 76832 39984 76832 0 vss
rlabel metal2 36344 73752 36344 73752 0 _000_
rlabel metal3 42672 75768 42672 75768 0 _001_
rlabel metal2 37576 73528 37576 73528 0 _002_
rlabel metal3 40376 75096 40376 75096 0 _003_
rlabel metal2 31080 74536 31080 74536 0 _004_
rlabel metal2 55608 75600 55608 75600 0 _005_
rlabel metal3 53592 75656 53592 75656 0 _006_
rlabel metal2 55272 75320 55272 75320 0 _007_
rlabel metal3 54824 75656 54824 75656 0 _008_
rlabel metal2 31864 71512 31864 71512 0 _009_
rlabel metal2 31192 75600 31192 75600 0 _010_
rlabel metal2 30520 74872 30520 74872 0 _011_
rlabel metal2 32032 74088 32032 74088 0 _012_
rlabel metal2 30856 75376 30856 75376 0 _013_
rlabel metal2 37016 72688 37016 72688 0 _014_
rlabel metal2 38920 73696 38920 73696 0 _015_
rlabel metal2 37520 71960 37520 71960 0 _016_
rlabel metal2 36680 73808 36680 73808 0 _017_
rlabel metal2 37576 75040 37576 75040 0 _018_
rlabel metal3 34944 74648 34944 74648 0 _019_
rlabel metal2 57400 74984 57400 74984 0 _020_
rlabel metal3 56952 73528 56952 73528 0 _021_
rlabel metal3 57008 73976 57008 73976 0 _022_
rlabel metal3 57288 74088 57288 74088 0 _023_
rlabel metal3 51240 73584 51240 73584 0 _024_
rlabel metal2 33208 76552 33208 76552 0 _025_
rlabel metal2 33096 74368 33096 74368 0 _026_
rlabel metal2 33208 75152 33208 75152 0 _027_
rlabel metal2 33544 73920 33544 73920 0 _028_
rlabel metal2 41608 72548 41608 72548 0 _029_
rlabel metal3 38276 73416 38276 73416 0 _030_
rlabel metal3 43512 74760 43512 74760 0 _031_
rlabel metal2 44296 73808 44296 73808 0 _032_
rlabel metal2 35560 74816 35560 74816 0 _033_
rlabel metal2 52920 73752 52920 73752 0 _034_
rlabel metal2 53872 73304 53872 73304 0 _035_
rlabel metal2 54320 75096 54320 75096 0 _036_
rlabel metal2 53984 74088 53984 74088 0 _037_
rlabel metal2 35784 76160 35784 76160 0 _038_
rlabel metal3 36736 74872 36736 74872 0 _039_
rlabel metal2 35616 75096 35616 75096 0 _040_
rlabel metal2 43624 71176 43624 71176 0 _041_
rlabel metal2 38584 74480 38584 74480 0 _042_
rlabel metal3 40600 71176 40600 71176 0 _043_
rlabel metal2 40488 74872 40488 74872 0 _044_
rlabel metal2 36792 72520 36792 72520 0 _045_
rlabel metal2 36456 75264 36456 75264 0 _046_
rlabel metal2 51912 71400 51912 71400 0 _047_
rlabel metal2 49224 71848 49224 71848 0 _048_
rlabel metal3 49336 73864 49336 73864 0 _049_
rlabel metal2 48776 74592 48776 74592 0 _050_
rlabel metal2 48608 74312 48608 74312 0 _051_
rlabel metal2 36176 70728 36176 70728 0 _052_
rlabel metal2 49448 75880 49448 75880 0 _053_
rlabel metal2 28952 74480 28952 74480 0 _054_
rlabel metal2 38696 75320 38696 75320 0 _055_
rlabel metal2 36904 74872 36904 74872 0 _056_
rlabel metal2 28616 74928 28616 74928 0 _057_
rlabel metal3 34776 74312 34776 74312 0 _058_
rlabel metal2 47208 75208 47208 75208 0 _059_
rlabel metal2 44184 75152 44184 75152 0 _060_
rlabel metal2 42168 74032 42168 74032 0 _061_
rlabel metal2 38136 72240 38136 72240 0 _062_
rlabel metal2 46312 72800 46312 72800 0 _063_
rlabel metal2 45640 73024 45640 73024 0 _064_
rlabel metal2 43960 71400 43960 71400 0 _065_
rlabel metal3 42000 73304 42000 73304 0 _066_
rlabel metal3 47040 73528 47040 73528 0 _067_
rlabel metal2 45864 73976 45864 73976 0 _068_
rlabel metal3 44352 72632 44352 72632 0 _069_
rlabel metal2 42840 71680 42840 71680 0 _070_
rlabel metal2 39816 71456 39816 71456 0 _071_
rlabel metal2 38472 73584 38472 73584 0 _072_
rlabel metal2 38584 70448 38584 70448 0 _073_
rlabel metal2 39816 72856 39816 72856 0 _074_
rlabel metal2 39032 72800 39032 72800 0 _075_
rlabel metal2 38304 74312 38304 74312 0 _076_
rlabel metal2 37464 72576 37464 72576 0 _077_
rlabel metal2 38472 72240 38472 72240 0 _078_
rlabel metal3 40600 71064 40600 71064 0 _079_
rlabel metal3 44240 71848 44240 71848 0 _080_
rlabel metal2 43008 73080 43008 73080 0 _081_
rlabel metal3 46984 72520 46984 72520 0 _082_
rlabel metal3 44968 73192 44968 73192 0 _083_
rlabel metal2 42280 73724 42280 73724 0 _084_
rlabel metal3 41832 74872 41832 74872 0 _085_
rlabel metal3 43568 75096 43568 75096 0 _086_
rlabel metal3 58240 75544 58240 75544 0 _087_
rlabel metal3 55608 75432 55608 75432 0 _088_
rlabel metal2 50120 74144 50120 74144 0 _089_
rlabel metal3 54712 73864 54712 73864 0 _090_
rlabel metal2 55552 72408 55552 72408 0 _091_
rlabel metal2 54824 75152 54824 75152 0 _092_
rlabel metal3 53312 74088 53312 74088 0 _093_
rlabel metal2 51128 73472 51128 73472 0 _094_
rlabel metal2 49896 72688 49896 72688 0 _095_
rlabel metal3 60368 74872 60368 74872 0 _096_
rlabel metal2 59528 73192 59528 73192 0 _097_
rlabel metal3 53984 72520 53984 72520 0 _098_
rlabel metal2 52472 72912 52472 72912 0 _099_
rlabel metal2 57064 72464 57064 72464 0 _100_
rlabel metal3 56504 70952 56504 70952 0 _101_
rlabel metal3 58464 71848 58464 71848 0 _102_
rlabel metal2 57288 71792 57288 71792 0 _103_
rlabel metal2 56504 71904 56504 71904 0 _104_
rlabel metal2 57064 74312 57064 74312 0 _105_
rlabel metal3 57344 73304 57344 73304 0 _106_
rlabel metal2 58072 72912 58072 72912 0 _107_
rlabel metal2 52080 73192 52080 73192 0 _108_
rlabel metal3 53536 72408 53536 72408 0 _109_
rlabel metal2 49672 72800 49672 72800 0 _110_
rlabel metal2 50904 72688 50904 72688 0 _111_
rlabel metal2 50120 72744 50120 72744 0 _112_
rlabel metal3 50120 73976 50120 73976 0 _113_
rlabel metal2 49784 73360 49784 73360 0 _114_
rlabel metal3 46704 74312 46704 74312 0 _115_
rlabel metal2 51016 71064 51016 71064 0 _116_
rlabel metal2 35504 71624 35504 71624 0 _117_
rlabel metal2 35504 72632 35504 72632 0 _118_
rlabel metal2 1792 76552 1792 76552 0 io_active
rlabel metal2 38584 77882 38584 77882 0 io_in[18]
rlabel metal2 42112 71064 42112 71064 0 io_in[19]
rlabel metal2 44800 69496 44800 69496 0 io_in[20]
rlabel metal2 47376 70392 47376 70392 0 io_in[21]
rlabel metal2 46648 71176 46648 71176 0 io_in[22]
rlabel metal2 49672 70392 49672 70392 0 io_in[23]
rlabel metal2 51184 70392 51184 70392 0 io_in[24]
rlabel metal2 54264 76384 54264 76384 0 io_in[25]
rlabel metal2 54768 69496 54768 69496 0 io_in[26]
rlabel metal2 60984 73640 60984 73640 0 io_in[27]
rlabel metal2 59640 72464 59640 72464 0 io_in[28]
rlabel metal2 61992 76832 61992 76832 0 io_in[29]
rlabel metal3 63896 76552 63896 76552 0 io_in[30]
rlabel metal2 65240 76440 65240 76440 0 io_in[31]
rlabel metal2 66808 77378 66808 77378 0 io_in[32]
rlabel metal2 69384 76720 69384 76720 0 io_in[33]
rlabel metal2 70840 77154 70840 77154 0 io_in[34]
rlabel metal2 72856 77154 72856 77154 0 io_in[35]
rlabel metal3 75992 75544 75992 75544 0 io_in[36]
rlabel metal2 77280 76552 77280 76552 0 io_in[37]
rlabel metal2 3808 76552 3808 76552 0 io_out[0]
rlabel metal2 23968 76552 23968 76552 0 io_out[10]
rlabel metal2 25984 76552 25984 76552 0 io_out[11]
rlabel metal3 28336 76328 28336 76328 0 io_out[12]
rlabel metal3 30296 76328 30296 76328 0 io_out[13]
rlabel metal2 31864 77770 31864 77770 0 io_out[14]
rlabel metal2 34776 76776 34776 76776 0 io_out[15]
rlabel metal2 36792 77056 36792 77056 0 io_out[16]
rlabel metal2 37912 77994 37912 77994 0 io_out[17]
rlabel metal2 11872 76552 11872 76552 0 io_out[4]
rlabel metal2 14056 77168 14056 77168 0 io_out[5]
rlabel metal2 16072 77168 16072 77168 0 io_out[6]
rlabel metal2 17920 76552 17920 76552 0 io_out[7]
rlabel metal2 19880 76608 19880 76608 0 io_out[8]
rlabel metal2 21952 76552 21952 76552 0 io_out[9]
rlabel metal2 3360 76328 3360 76328 0 net1
rlabel via2 56280 73192 56280 73192 0 net10
rlabel metal2 7112 76664 7112 76664 0 net100
rlabel metal2 9128 76664 9128 76664 0 net101
rlabel metal2 11144 76664 11144 76664 0 net102
rlabel metal2 13160 75544 13160 75544 0 net103
rlabel metal2 15176 75544 15176 75544 0 net104
rlabel metal2 17192 75544 17192 75544 0 net105
rlabel metal2 19208 75544 19208 75544 0 net106
rlabel metal3 21448 75544 21448 75544 0 net107
rlabel metal2 23240 75544 23240 75544 0 net108
rlabel metal2 25256 75544 25256 75544 0 net109
rlabel metal2 56616 73192 56616 73192 0 net11
rlabel metal2 27272 75544 27272 75544 0 net110
rlabel metal2 28728 76160 28728 76160 0 net111
rlabel metal2 31416 74088 31416 74088 0 net112
rlabel metal2 32760 73808 32760 73808 0 net113
rlabel metal2 34832 72408 34832 72408 0 net114
rlabel metal2 37016 72128 37016 72128 0 net115
rlabel metal3 37856 72408 37856 72408 0 net116
rlabel metal2 41104 76664 41104 76664 0 net117
rlabel metal2 46648 73752 46648 73752 0 net118
rlabel metal2 45584 71960 45584 71960 0 net119
rlabel metal2 54936 72688 54936 72688 0 net12
rlabel metal3 47936 74088 47936 74088 0 net120
rlabel metal2 49112 73164 49112 73164 0 net121
rlabel metal2 52360 72800 52360 72800 0 net122
rlabel metal3 56952 76664 56952 76664 0 net123
rlabel metal2 59864 73752 59864 73752 0 net124
rlabel metal3 58856 73864 58856 73864 0 net125
rlabel metal2 60424 73640 60424 73640 0 net126
rlabel metal2 61432 77378 61432 77378 0 net127
rlabel metal2 63784 76440 63784 76440 0 net128
rlabel metal2 65576 75544 65576 75544 0 net129
rlabel metal2 55384 73696 55384 73696 0 net13
rlabel metal2 67704 76104 67704 76104 0 net130
rlabel metal3 69776 75432 69776 75432 0 net131
rlabel metal2 71624 75544 71624 75544 0 net132
rlabel metal3 73752 75544 73752 75544 0 net133
rlabel metal2 75768 75320 75768 75320 0 net134
rlabel metal2 78008 76440 78008 76440 0 net135
rlabel metal2 5768 76664 5768 76664 0 net136
rlabel metal2 7784 76664 7784 76664 0 net137
rlabel metal2 9800 76664 9800 76664 0 net138
rlabel metal4 39928 75656 39928 75656 0 net139
rlabel metal2 59192 75712 59192 75712 0 net14
rlabel metal3 38108 75432 38108 75432 0 net140
rlabel metal2 47376 73864 47376 73864 0 net141
rlabel metal2 47040 72408 47040 72408 0 net142
rlabel metal2 48216 73164 48216 73164 0 net143
rlabel metal2 50288 70840 50288 70840 0 net144
rlabel metal2 59864 76496 59864 76496 0 net145
rlabel metal2 60592 75544 60592 75544 0 net146
rlabel metal2 61768 75376 61768 75376 0 net147
rlabel metal2 58072 77322 58072 77322 0 net148
rlabel metal2 62216 75152 62216 75152 0 net149
rlabel metal2 55272 71232 55272 71232 0 net15
rlabel metal2 62104 77154 62104 77154 0 net150
rlabel metal2 64288 75544 64288 75544 0 net151
rlabel metal2 66360 76440 66360 76440 0 net152
rlabel metal3 69048 76664 69048 76664 0 net153
rlabel metal3 70448 75544 70448 75544 0 net154
rlabel metal2 72296 75544 72296 75544 0 net155
rlabel metal2 74312 75096 74312 75096 0 net156
rlabel metal2 76440 76104 76440 76104 0 net157
rlabel metal2 78176 75096 78176 75096 0 net158
rlabel metal2 73080 1134 73080 1134 0 net159
rlabel metal3 54852 70392 54852 70392 0 net16
rlabel metal2 73304 854 73304 854 0 net160
rlabel metal2 73528 2590 73528 2590 0 net161
rlabel metal2 30296 2030 30296 2030 0 net162
rlabel metal2 30968 2030 30968 2030 0 net163
rlabel metal2 31640 2030 31640 2030 0 net164
rlabel metal2 32312 2030 32312 2030 0 net165
rlabel metal2 32984 2030 32984 2030 0 net166
rlabel metal2 33656 2030 33656 2030 0 net167
rlabel metal2 34328 2030 34328 2030 0 net168
rlabel metal2 35000 2030 35000 2030 0 net169
rlabel metal2 53200 71064 53200 71064 0 net17
rlabel metal2 35672 2030 35672 2030 0 net170
rlabel metal2 36344 2030 36344 2030 0 net171
rlabel metal2 37016 2030 37016 2030 0 net172
rlabel metal2 37688 2030 37688 2030 0 net173
rlabel metal2 38360 2030 38360 2030 0 net174
rlabel metal2 39032 2030 39032 2030 0 net175
rlabel metal2 39704 2030 39704 2030 0 net176
rlabel metal2 40376 2030 40376 2030 0 net177
rlabel metal2 41048 1246 41048 1246 0 net178
rlabel metal2 41720 1134 41720 1134 0 net179
rlabel metal2 70952 77056 70952 77056 0 net18
rlabel metal2 42392 1302 42392 1302 0 net180
rlabel metal2 43064 1190 43064 1190 0 net181
rlabel metal2 43736 1246 43736 1246 0 net182
rlabel metal2 44408 1134 44408 1134 0 net183
rlabel metal2 45080 1134 45080 1134 0 net184
rlabel metal2 45752 1246 45752 1246 0 net185
rlabel metal2 46424 1134 46424 1134 0 net186
rlabel metal2 47096 1246 47096 1246 0 net187
rlabel metal2 47768 1134 47768 1134 0 net188
rlabel metal2 48440 1134 48440 1134 0 net189
rlabel metal3 51128 71008 51128 71008 0 net19
rlabel metal2 49112 1246 49112 1246 0 net190
rlabel metal2 49784 1134 49784 1134 0 net191
rlabel metal2 50456 1246 50456 1246 0 net192
rlabel metal2 51128 1134 51128 1134 0 net193
rlabel metal2 51800 1134 51800 1134 0 net194
rlabel metal2 52472 1246 52472 1246 0 net195
rlabel metal2 53144 1134 53144 1134 0 net196
rlabel metal2 53816 1246 53816 1246 0 net197
rlabel metal2 36008 74816 36008 74816 0 net2
rlabel metal2 75096 75712 75096 75712 0 net20
rlabel metal2 62552 75152 62552 75152 0 net21
rlabel metal2 6552 77000 6552 77000 0 net22
rlabel metal2 29288 75992 29288 75992 0 net23
rlabel metal2 27272 76496 27272 76496 0 net24
rlabel metal2 28280 75992 28280 75992 0 net25
rlabel metal2 29400 75152 29400 75152 0 net26
rlabel metal2 29512 75936 29512 75936 0 net27
rlabel metal3 33376 75544 33376 75544 0 net28
rlabel metal2 34664 75768 34664 75768 0 net29
rlabel metal2 39592 69944 39592 69944 0 net3
rlabel metal2 35448 73752 35448 73752 0 net30
rlabel metal2 13832 73584 13832 73584 0 net31
rlabel metal2 15848 73976 15848 73976 0 net32
rlabel metal2 31304 75264 31304 75264 0 net33
rlabel metal2 20216 75376 20216 75376 0 net34
rlabel metal2 21000 76328 21000 76328 0 net35
rlabel metal2 24024 75936 24024 75936 0 net36
rlabel metal2 54488 1134 54488 1134 0 net37
rlabel metal2 55160 1246 55160 1246 0 net38
rlabel metal2 55832 1134 55832 1134 0 net39
rlabel metal2 43456 70168 43456 70168 0 net4
rlabel metal2 56504 1134 56504 1134 0 net40
rlabel metal2 57176 1246 57176 1246 0 net41
rlabel metal2 57848 1134 57848 1134 0 net42
rlabel metal2 58520 1134 58520 1134 0 net43
rlabel metal2 59192 1246 59192 1246 0 net44
rlabel metal2 59864 1134 59864 1134 0 net45
rlabel metal2 60536 1246 60536 1246 0 net46
rlabel metal2 61208 2030 61208 2030 0 net47
rlabel metal2 61880 1246 61880 1246 0 net48
rlabel metal2 62552 1246 62552 1246 0 net49
rlabel metal2 44016 72408 44016 72408 0 net5
rlabel metal2 63224 2030 63224 2030 0 net50
rlabel metal2 63896 1246 63896 1246 0 net51
rlabel metal2 64568 2030 64568 2030 0 net52
rlabel metal2 65240 1246 65240 1246 0 net53
rlabel metal2 65912 1246 65912 1246 0 net54
rlabel metal2 66584 2030 66584 2030 0 net55
rlabel metal2 67256 1246 67256 1246 0 net56
rlabel metal2 67928 2030 67928 2030 0 net57
rlabel metal2 68600 1246 68600 1246 0 net58
rlabel metal2 69272 1246 69272 1246 0 net59
rlabel metal2 46760 75936 46760 75936 0 net6
rlabel metal2 69944 2030 69944 2030 0 net60
rlabel metal2 70616 1246 70616 1246 0 net61
rlabel metal2 71288 2030 71288 2030 0 net62
rlabel metal2 71960 1246 71960 1246 0 net63
rlabel metal2 72632 1246 72632 1246 0 net64
rlabel metal2 6776 2030 6776 2030 0 net65
rlabel metal2 8120 2030 8120 2030 0 net66
rlabel metal2 9016 2030 9016 2030 0 net67
rlabel metal2 9912 2030 9912 2030 0 net68
rlabel metal2 10808 2030 10808 2030 0 net69
rlabel metal3 47992 73304 47992 73304 0 net7
rlabel metal2 11704 2030 11704 2030 0 net70
rlabel metal2 12376 2030 12376 2030 0 net71
rlabel metal2 13048 2030 13048 2030 0 net72
rlabel metal2 13720 2030 13720 2030 0 net73
rlabel metal2 14392 2030 14392 2030 0 net74
rlabel metal2 15064 2030 15064 2030 0 net75
rlabel metal2 15736 2030 15736 2030 0 net76
rlabel metal2 16408 2030 16408 2030 0 net77
rlabel metal2 17080 2030 17080 2030 0 net78
rlabel metal2 17752 2030 17752 2030 0 net79
rlabel metal3 50708 73528 50708 73528 0 net8
rlabel metal2 18424 2030 18424 2030 0 net80
rlabel metal2 19096 2030 19096 2030 0 net81
rlabel metal2 19768 1190 19768 1190 0 net82
rlabel metal2 20440 2030 20440 2030 0 net83
rlabel metal2 21112 2030 21112 2030 0 net84
rlabel metal2 21784 2030 21784 2030 0 net85
rlabel metal2 22456 2030 22456 2030 0 net86
rlabel metal2 23128 2030 23128 2030 0 net87
rlabel metal2 23800 2030 23800 2030 0 net88
rlabel metal2 24472 2030 24472 2030 0 net89
rlabel metal2 47712 71960 47712 71960 0 net9
rlabel metal2 25144 2030 25144 2030 0 net90
rlabel metal2 25816 2030 25816 2030 0 net91
rlabel metal2 26488 2030 26488 2030 0 net92
rlabel metal2 27160 2030 27160 2030 0 net93
rlabel metal2 27832 2030 27832 2030 0 net94
rlabel metal2 28504 2030 28504 2030 0 net95
rlabel metal2 29176 2030 29176 2030 0 net96
rlabel metal2 29848 2030 29848 2030 0 net97
rlabel metal2 3080 75544 3080 75544 0 net98
rlabel metal2 5096 75544 5096 75544 0 net99
<< properties >>
string FIXED_BBOX 0 0 80000 80000
<< end >>
